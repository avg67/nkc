--
--Written by GowinSynthesis
--Tool Version "V1.9.10.03 (64-bit)"
--Mon Apr  7 19:25:26 2025

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.10.03_x64/IDE/ipcore/FIFO_HS/data/fifo_hs.v"
--file1 "\C:/Gowin/Gowin_V1.9.10.03_x64/IDE/ipcore/FIFO_HS/data/fifo_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
Afsfzdw9aSU9h2ZGKzNqTBSyu99yiiFyXVKq0nRTjlB/YwcHLVCXqwGbKul3O5fMdBQCYdDchULx
k2OJThfCEM96QX6JP9JtQou/hjjZ3KOKwt2sXt0icK5FrHU8i5pOvLSDoz/NVN/xZXAHDuXF+5Am
E3jXXaLR0t/IjjQInhZ7NNzKuLsvzJTe+dQOjiDkIJK3ERR+pN47ffpG5TQW4oBRXhDiQuhN48ZS
cgA+KducMFOSwjWoOk/DoQoUilD44ybDe467CUkfYhkbwQOBz7CvXiyzhou9tJk3hWuLqK0l2rkC
ypSypIj7e/Aj33WRk1Bs0dgPjD7zRccDIQSdcQ==

`protect encoding=(enctype="base64", line_length=76, bytes=21888)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
o/Liqf6xctI1MrzLCcEtXGRW6n3C1TdZYdfHwHBaE4fWJjQTM79wXYYRTj7DP47LaP+IY4wfByi3
C+Lu+z7qKr9YIr27bFf4SeEmS01gWUagUNSSMk5Q5tvKneeHxvSNez30VIUBwNo2qoexGEFPc+Hg
zEo70MJ33UWEk9EHwM6cbHxxt90JV/e8jMNw4UdOy0rj8bY+NjwfxY6WFMf3HI9Kipq/WP3ORwkV
TBpdZc7zm5q0r3wpLbnVMvyELA5VRCyYeFJ3LGR8V4kZa/9U+PoyLunxpnK6my5v43z5TPnJoHoA
ymbI5VfLStKKjCD+yY52Zk+1u6bdCmF2W9mcHYlVQ6Ny25YkaPytnaRa1wBt7Neb3EoG8bEggbgx
JZuSiI7hwiHg+Fr9QW2mCFrAB/wwP06ELfaHBi7+OASCY5cV0zEV5oHJZZvbFZVtblHvLHp2F1bi
sPo3A5Nz2ImYmBf6+UO3b+UPhgL7GoKP0pLuaj44Htd19m1EcM7VR5w029wu1a33gMZzEBeeBySH
KHod85q6bnjciH90Z+JTEBWOzajeiSq0eNyechWMdRV/gDo3sFduffIhGLD8HlxtkbDayKwtYGMA
is8FdLRytiZoyHXr5jMphOkRqlfPmgwy4E9VaexU0ouXeTtGs9tp4dgWyMUvwx3JcqkByRaf0O35
8MNU12ylstiVhAbzDxu+3c5e9exY97geX/AhL45cJKx4brBeDSE4/MHoX2up7esHU3Qa625twoo6
o6tMYqe5dmxrkZ5xg0ukLevzg3dbdPLljdqsq/Itd9L+cFFkffOld9FWpo+FWh1KouoStgqO/NGI
eSAPXWG4f1foKYBhHPvz49RDy3L+JAKYCZm3TpSUophOxUnlBYFGVW1pKKqCXACcLAeDtkED2R5O
HLVKoZiXVHuI8Bb4a+5FwTYa+RhV6J8Ect92E0g3n7xu8kR9ror1VL2UQ4w9zNNhpBsvg+3QFSYA
R35ZZvuik3M5gH/qofw0N/XSFs1dXOMrOsN2nzGZ42NIpAR3vXRYSOdK3lm4V8nwUXhHeGk/UbMo
La+mmDz6JuyDJRyQ9OVlLTq201epCf/UL2js98rgFJq8utdXKpaEKvs6UtTxx74Y44mvhCIhrgVE
KrV5VMf4Qq5+DyTyb3PS+TkyDsedL+e0Z6WnFj6DiQPOg/RBBRqz8Ifp8MNGp1LO0R9XYcepKpIq
LMyZKr/OQ6oErKWixEx5tlR6iQ5ByKt5ellkqKlrX3hRbOdOO/QkJ4nwKqL73Wr93V8768w6nsZg
t8EY/WbjgkER8c8R3nP7RXIO7qe8jVKFDLaEJTIcWdQfPpAT+ofEUm7M0DK2fSxxu+oq/F+OU817
ITn7Xv1G30khA7v6Krm8/AqjC8lyT2wGz/auaw1lHSOazjjT0RFaOrDwbJTK1vEw43abVZjyIFAv
Qljmk1MZJNy35GFLt5XMAGrUIVZ6eM5d5Z1q8djSB1bFixm5CyyoFZdNyAzpQvkN6Or7GVehQU/x
y54TVmKsOx9zfLrgOqch0pn+CdQzaLcgFzcn9LHNbX2JHmuGTso/gq8Y/OO3WQd2iReAyEgy2+om
u55hTcket7XQKIhwzvDssuQlurDhVz5uwqX3sB2JSZwhvCTdEwH6sE2Zurv+YvCLuiU6vwmy0NcK
yky5r6FfTPfWmPvfn4vNrKH4ei+QTjv1o/Wm0pYXnRpjpcEWKTM/OuoNAIZER44rmNY9YqDCD3jN
fkA3vXWw9iLB2Kr8L5s7FqWxm9wKeTdiFzqm37tIgeZ9uMmIw1993MiVlCWQUDRgedDd6YN527WC
pHLT4v1pwpa6SU1unWxxUxkL9s9KMtw6ufwh1ZYilQNpjuMoRHV6pfBJQRLdGsVnuVu2x4K6lxlF
rka65D6mOLFmWG0me+7JY2DoD6BoXNV9YGbuVgavkXUpIpeEYc7xk0YNJWDIlotB9CNTNdh1LjsP
NaV3ZPKt9k5ZphSwptYE9TASbowggy/YsUw9w7xP6R8Xs8sI7RbIQ8Mv1VVneK02A44CKlsezRva
BM/mVshNggqPg/yZcSlkpGDYNW6vnjAFURAbRnhk5ICOguaJKjjq0YFOPZWWnyidOXLyrr+4PI6E
H7UfeRAE+dBXatr2xT3+nQ3oeyLgJHNLMO03wTRALQuDUxLHJQZCfwSExy40sN3QOYmND3KzsV5t
7Lmo+T7CogUCq9zC0TXz4meqDkZNOoLI7JF3hn+0Vg45NyKZahecwcFXH2Vh0akw4xtosagVWJRc
xaxfZ4TxLanLpvmUbnEU5gPxlWc+M/DW2VY+vMkpYV6uzn5dSizSR2J6WjhoEFwrLGzmaMu+cA1F
FXOaes6syGlcovIP3LvB7XnHGz3kP4DNuq05PhyGvsKlHDHWlDJg7tl+dH3rKaN4vdmksanfTerD
ygR2grlg2oXz6Ni7VBMcG6/BdqZ2cxmeXJGQwSCyk/OetsV6Eb44mSIKzZGX4sz29xkSWU0lB/im
09WlPIKe6EGkx+hPUtOgxOFgCKwaomwfBvn8vhiSPweozIebHBmw9tJ7Jujf29mRvyOaFyS3GMXI
qkd00uWiPizv4pjl7m8n5E/F54cc3v5RNC3pOKqlSnvQmwi18L7/PDvUz24gwv/m7UFOM3qHtekw
PnJRIue52F64cwe+hrnjefwtGpW1Fy8//WCTe+EW4ax5HaI9tt5XZf/uyd8LGLhJwDIKhrUBzb79
uZMrpjVW8YtxpAHJ3WycyBn5WfxsBVWayVhSqZRf1MunZGcEmwvNIn8jNy9uPaG10H2FYpv9cxgz
6zzhByQtNGENRgDkUXe0ggxWuXQ2pug41PFWiSYGYkdL6brRdMcJ8vUKpZkqSghCZuIsHOxPbNdQ
FsngeXLr+dcidaC7oMaahUzj/WcoYmXQUXXho8Pk6yR5c20974e0XYOIHHCD2V0KrM2CPY2n18MA
06EcR4MFeeDdgddB4hMIH11aMAVYy/WisDW9ZfZxk8SOg3PW5y82wtrRAtOoEjXMFI51yZiWwW0C
qcIgUYlzHRn4c4lYiN0r0sbwO1MMeIORdZDLX0njb7/lQr0+127QsgNkxw8UNIkvTcys3drG6vhK
CLaHiloOpyGgr81z+UJA0IGl3eR5YbJnqSC0/0FTRH/44WHC+/kcyqyxBC0NJipwUUmD4BdLRDt/
7KOID0QP8kR80uNvvMTZpNrRtUsanBIRdPD5rQLnCrgR4i2OI/pBH5iOWWf5AarKXZYnaufFdWKm
aFObIkuONAQ6oXlGYLdXMyMbM+UYK9bgUmDNsOcXP4ibRFFf3jCGMAB/c4p3ye46M6VOJMACQpaw
7Pese47JyZK/d5RXKGp4Sc5vQfNnJtrDzx3J0iZB0yc7QgEzIF62G0tOTx2dIBARMn/6o3KIilxA
I2krqDna/TuJ/UCUNYtG3nha3CJc0YOLElypZ8lwN7+DzZL0vbQnQpSMuhu13tqXKoAO2KcskU5O
BEuNr67YlV0BpBhtAMyZvGB38uxN/oPoPGlDfprg+NW5YwbSr/UMAdqwSSizVEEsBrJeEOyDhgP9
OMC7APKUFduhU2KnyYbEpJ+Yt2Ea1V0CSlcAxlomZEW6ON/m/BvfxNU5ioqo3NQ85/Ca4EzpnUN5
9pkXJls6rgiN73RNTo14Rw1QmcZNF7DHJxco4CuqFvOZFwhEGRS/Q23ej+kU6cYT9roZ2yfT4z42
eXPYGRgx0z5/Yl4XYDhW6hP5uoF5uc/sYh6H17fagsdEbBQXsZ6xwz9QxhYj6WxV4fdJ/8heJGuI
nZPN0K6RiKPLGfX80oIgEXF7rYHy7XHngJ8dRpJY4FLD25LMpTc90AjaLZ2FeJwBV48tuAQFKu8o
l2ASYzYdLWP+xU4Q9I+/zTXYU29OUh2U8AGtZ8fw/2MnfaVaqeSJUWK9ijh+n1U1efXEi4vPhgaU
YY1e+NbWwgE2sV09ZGkgbZueT3iOSz/qOH6D1NNvD96RDFbuUbNfoQkjinJ+5TVie6gHyQAxww8w
/CGX+1YGy7PE8FbvfiA/WVxkbOZK3bINW4Lm+EshqvReehBwLymyIQt2BUCID+gFD1vHRAjnFfDG
YIhUVH3o2MAkP79VOHm7ntE1KNpVsctvHxOks1yi1+31Dwbsj7JtM6PwcbgmfBOE6qDt7yw017b/
BhC2VDaIAwfUS4AaIzQy4YclA1JAk17U7VKcsBZh0oFYcvxlkirROhUaPm6EiSNgMRGRU2BXJKNY
GkRatbEeR7lET851DHQhKOXoWYrodzb3wfrSTVivvZfMHZT849WLh8mFBKId23UCM+Opxn8q6qIu
o/NCX3VODWZCD49KbrjU/ThpfloODZ8EOFRIOdk5Fdk7McTvWsNRxDz6a+IyYnWPaxxRbeho8A/3
vfosJ/PUHrlO9929RV/gWuchbBIczMJPA5po1H1G4E/2tsdnZ0XTxnH+loytl1gdkP+nqdSd81dS
+/AjeF4lcYZr2zWywsCYYX0P3O1MAuxqcxWXeui5uOvtRxudi2HkBDsNnzrZymbU1IZRLQYPrV1u
bb9lIV9O9bQ3hXlDQtY38jQQN4dQ7CUuCO/f07eAXlndFpdZQrVaIprNk348Xg7Tm3izKbyCo1wU
kX7HaoNPZDlqE9E7PLdGKAAjHhtAE02tCzYdsfEkoh+EMghP1wMIFK6P+NKymJdyqD9RhiOWGKSt
Nny+VQFz1O2gWkGGhnDkxpDmL0t2jbTpvlgS6jsZj6v209K5MMzw9l4Kk+4SbLYVj46j/9FfaYJZ
3c4uBQX0Xdksk5e0FBNJCoaPw/000+uYXz/lRo+hwK/+4ygofVozR3daq/9XJgzJRER/KHpoB5bH
Q49h/jz8VMDLhxLs+nTUtXslumSRxQgfQqqoFW+Pi9YeNZkw0YmVmsQ89SiZ0qO5pCIvKpjSipnx
H9c1HxytIodvMRRbWBTvG1nttHX6ZuP2cI9hdWYDcJqhBo60CqxSr2PNFRonkKEiffyap09xsbSY
YmjW9ggVBXvMeMvdhDnkv7wWMoNmAzA94SrDEug+8UzlVmH8KI3/WKsJUl49yvTJUsVl/no0gMcF
h8uQZA7j3JB2r+kP2Mu/CQ5YEt2q00mUvmqNpZgVfnfy089gTQ2MC26JDyMrg1NDT9h9kaAQfBAz
03nmCl6ttbW/YPP5rkMt0LmdZBpVmfLdWyH3A3dWo/Cvsm7uG2qNhINMd96rTTeAcear5hzpUoce
7rVFfooz+ZUpujiBrjY2H3rbWzKbUrsjivRrS/j8MB2BMlzBB+toxn90ta3YpIo2eWKm8DKP5D32
Sd533poU/Of0uzGbt96gHp9jQitN8zBp6OmALkIPMyxTRI0mpR1LU58mJ2Dzy4Tt4JJx3H5KjJEi
905CtnlF4NqC5mYDNRKhM6YEePD7KIwmjkdi6oYOCwe4QmgizR8JsX8zyGLaNGhgZIMFRsN3j+lA
zMEy0uQHesOlYAMSnJ1/XpV1xfqM3SmPA1XdCvBLx4JeUvYR4FEeHdyRgL6YY7vVM81nH26Z9ikZ
SFJxRU/tiG1KtJ29QUBKJFBWk08c/9SUwdJmeE4vemJJNSIO1F8e9SSbksvRL6KNIs4jcAQsquIJ
XulkkF9rdHPnz3byOEG661HyKy/l3HaOCOphJsilPEAJyQ7jWGKrSOfkQg//tZsMs2xBJF89QtZF
orTQ7Or2mEzLPbXDiVmljHLgF/jru7MZFF4tSSGbReuhYZyLURtTnA1T3U5RT/n+rpnAD9cnTewn
RH7H8VjssDu+L6pPnUAj2YpjultpowB4oM/1DCkxa1JYyzq6yCdnuUlnnj6xyyN+epn5lH3gjx7H
gtvznvMrDYmZaP3PqZNkySdhLS6EAnvYpIQyPdZyoMIYtb9PaEs4BGFQRXfJ95OMsngFmKR8mkyb
4q+vULLTBDRipMR3Hk+Ik7LYZ9BOrifozU5yiiqGFIse7q+WEN+cFsDZS0sbDv2+z32Cav6yn1a7
J7t3UjMMzrhNbZy2Wi/ixhSup+cmj9gZJkaG4GpnMcbviLBfnWQHr3L1IdHVJdbNbdcQ1O/UYXdz
9mYd1/6Bp7PqQGzUpjhrjzGhidO2ezvUdUSyWRW1sUgv+rEQVE9Klcm39U0/S8czqn1h905yy57z
p//Aq1e6URJ3gbbWCmqTaugFrU0/gfd96FBEKm5TJJpc7gS5eAHKV+3SpGKExSIdsyjXdMP6+AeN
9O6QJk6aSdyhsGQ+f2iBJrDJ4vaCN0HjFoRX4MpU9h3IJVHgaEtP/YYIpvCF5nC6Vuxd3NjJCPBp
rxC38PLBBPCxVFlDeJnKEo4DFFSIt7FE8ja/dgyEuHhDChBQW65DaJsSUXX9GQSN4yrxD3qhy4HT
D0lruZUgPqzIW4iAf49ez4tR0DzGSkTM019PPJQ0DEziZIjo8CUxq2ygRmGcENeW/Wkn/dKUeswj
VlJ0D1SBTC9ZdJtPn3oi61VFuIoWx2nOv1QhiQIFbhJsfH9mC247dneT2Pf1fDXutVnzyscUeDoY
06xaKaLKM+d/lsVxXhkVG2eHT3tYhnM+ri+G4xtbaLCukfBU6eYk7Qq3nqDDjJX/GgjXxgJx+42e
6hKT784XcbryaphpwmbmTTIOOHWjKmTNpH2IstXKzWTP/s3zy1tiDtAphwTbs7PWqJXqLtFoxKI8
V2F1EFy6+a/Z6aBgmGsIh7X67/5Ic5QbG1x835UKLYvgHBoLEdEhkdYNhulAK83ydHenhumsDj5x
tCqvpvQBiaAZCwn1uMRXh0BA1OhPb/MFKafKMizCQtgWlnc/GPS5ltm0W4e2Ny7/yeGNJzqxllMr
B6z5s+xcX5R+/e//04YvWyXazIXuf5hrOB6ypA7In5xJ9YWOF6LurFLLBARyXvIdIpF1woplqD1D
a4AA0QE93SEIa4Te/snM5Kf8owqCJsMpZKG2OAz4z/f1P2aUrbAeUuglTY8MzGCMoN2sfDalfQZA
vuPQ/dEDHvhAh2ol90HkJsHz0sltQ9Xkj+UNOkHEM8YP/LPHbeIqTKyudXEfjPlsgLQsH0GXP9u4
Vp6d2cuQq1KNOZ8c8n8SN4YzhCbfnWeoHmhfQ1BuGGLxo/oVuZpqmIxzQp/eUkSN0Mhx2ZU1M8E0
1vp3mVoRp/pG3izGWUdheuRWedz5ei3PSIN3ZHKZ4QcIYFzeLPyGziQRJoz7OIjfXjEeen3TQVbS
lT9IvfPw/3ubo2c0naozCF1Fpv/19WmzaP+hyBDxiltDnfL4T6mfEkjnthE8eT9jL0iWgpwTGQ7j
a+QzWwcqp5YD789+PSn4cgUYiaLk9tXYS6sWzRV1zMjoIcCf1SBbgr03eYtoV4o3dEDhKuTacvN+
Ccx9K6vzbE345izIZc+wRvhaQtmfGQb1TUZPG+2zahXd+M4Qy50AcWsFK+ft8JtvM56y3w5flAMb
6TyMsOAm1neDoNyWSBlDQ7gjN2SurJqplU8toLZEmbNEz3WsV7lFBs8MwFPBu1lPCrPkzkXAAHiq
3BqO7fjkEQ9nEhoMC5VOroDRkIEIhAxADhrLhvTXTeg6CEKTd8ZRwyGBoNjhUJ3flz939ZDKUqq+
hKx9JVM17XTT9NAD/yzcRamYwWq3eOjTx4xbA12w6EZZDVj7TLagxFI92u/DpzU+iZFO/D5heCUx
4rB0cob1Bh0xX5Q/qXM1YSGPOPw1yq5w0uNyur9lkvso02MbEiGZybTTGBvjN/96L6+iwvAUNDkM
jA2VIlTf8Dr/QQwIj0o7osE/xDQ2lqOnl0EvWxUkLUd9hAKmJ49yP+ZvMiWQLquRQ5niiFtCl290
KtzVkLSliGX6m5V5AdDK+y5V1DQjrlcC6sAB1Nst3XNUy5kF6Pi/geWJdoSBU3bOvpD2sy75pYfo
q0sekh/mxNOn8GjX1/J+lR1iGX31egbaYT+w0/RxKauPx7vT6BiaNwyj00bMckMsJ2lpE3JamFUo
46AcmhCpdgphZXlIqnfVTKiJhWU/imhEievxIFQYmgjrKvF5JhN16vwuhpUr4Rxq7gZas0SfHT6q
WZ+TB24fi+YKlF2onBvhykTEgjRdtH3bf7p1TrRvY+vLlH3tt5G1mrZC/xIiJ6ze3F3Quyvehqs/
aBr5UV+GT4k0mqg/VotK9KXGf6e4g+O//bB1hYy1mn7FwCN267s48Wy1cGNkiemiPjh9RXHVZmbv
fNEo2vfNnSs9R3bpx/nqu2sKBtgk/rG6o9ijCIONvvD5Mp1aLFTA9Xo9S8NSymL5vksELbTN1UMM
Gswkhmz7IB7GiDKaDi/sDajgEKiBlG9lVcN36lnlgtjmMXwC7UXF4Wo9/MYhtDUeFZF8J2/8/KoI
Kb0VWUMY5NNPmmutBKEpyyER0hiWfgFxNIeKZaQhSg3iptsm5KXGyPr5pVTH0LZBRnb8ImjEUgbo
NFkahCz1Fpe2mmc74EI1bpcmWeb3JBWhT9a9AklGQSdJOAsv4wrW0uMGiHv0SZQ2UyTDwCS/9ocB
GIrWf9FIat0kg3zhXkXcku2f9kh1fJCRDVKRAJ4ftyx80srIrUrIqKJdlHh/MrpbMVKRCqUDFJrN
vcLe9Xclcxj7EfxylfwZAIYJU3pRJhMbEbvbuvjp+CtWI8MRvkpYO4F4fR6uBmabICSmGMa0X59F
OBQDWKGrpdPa+9X/ai1V0ql1w1U5KBhzQhytAoCUpaYIMLy0Zz6dcoOEqZb7DEBYUVddYaNae2Mi
W/887ViLLOtVXNEvl5XCwsIEf3PRZmv8d0T3DC8TpMg3IucUFdSbYaMnXwhziUoAgG3A6vFc15dQ
B34IiFPj+BHUrWOnVSIpgkUhKq+/4a9GWZFUelS1ioiDATzt3SxdumMI8D/uX0HBWzjIg6vQUWIk
Y6ppmbYBEeOzEfPf8aZnN56Li6UGBIRwl681gTkJNTN6ErI56zHpCe3rAodwfF3ka6jJrG/3WiRE
lReNDdPW8VFulW0K1hfPzlRyk8p1ev7bCE+m/MzJCLelWYbfU88keSpFeN3nhCG/GOQNswvXhJfb
wg4ivPcspowMqTS5US3nCMUIcUrG4JDwJuewKDuwgLbysQHZ1+m4qxtWY+MHEUWHG4EG89kfTbKN
qiZuE/NxJEgO9lHMjAbWbhmk7wP0q93X925k4voxpKEhPhMhvaE5pWeKUyWr4IVfEdEUYyLWH8b3
0VZaQfTsCFtedQGbY7Is7BImv+Tib44+mi1BoYiGvGVtHRmpu0Vg9Vbpp5t4wBUT1Hg6FbUCF3bV
t22CDgsOfsg6iebuv4IM9/C45+65t6J80LO2Ed5nNxLGNxWKPh9u6+ShkQogy5c9LPOLu7TjMwBU
2yxaeZnst2fxhHdv7ohl67nkEM4zeoVWYE96zkTqgFUwsQTg8YXqVvGg1VNHNX2N2bQGWkhv3Fed
87kHZ5S7MjbWNJ73a1ar/UGiEP/ElhlXcPRhl4viZVyX48OgqKbGET6MMgYL/McvIFhmD1vnJMPP
qrVDo3/R4mYGprI8xRJDu63nfYLocJoZh3lO20Noror2j5XSEfmMDfAtqI/Lst5C1HOVX1LPkxQE
05B2uf0hcCYeWA5ZkLqEASziFFxqm2fVVS/6JpJxim/FsuIuP2cYJtw4dj4XfcgoR6bt0IUav7B0
F+W1KMnFvS8QK8Zsv5q6Y9Ppu8e8d8DXEQLpziGlQEDYJfScnENYQRHNz8Y23oqRQwe5VdIhmZk3
v7WI5WKe0grgB9VJ+3mLifj5MPxO7/AoyiMKW1T9d5QVi4DH9I5rZS0HobMfUYWq9MZm40wVzpet
k+crSibAFreCFSs2efQIdhvWyLtcihk0t2tHxiLSjK8pRj9Qsz8pM5dPYsHcXY7GpuXLQJXLqSzV
hxRhlVhlWSo0BenxOPS/suXcZxAiPlSbBxnVUJHcpY5siI1MwB/DyPPDJ00EsgSqIGsWJZ8zDRps
q7Xr5tQE1i8+j0nZ+NgAohC4kqsUdOU5E586xyF3NNmACTBfNEJFQ0ZGfJtmyO66enMAMD0dEvX2
MR31jTptFo8LICyJUa90sFoHfpCs4LcBcmfY5Ho2zwDmCHSmp9hC76YbcjHAWQv37BhFwOFe7FhK
g3IwqsslONiNmzt3RblZClGhlc5ERz2XW4oMFm5P7BVg8EXmBaQTtZsbXsnLjKbZILx5WWKTzb6Y
7y8n8BBfbmFONmJZHYqW/X916WjWfrC6Z+T1Mnua5NNbuYHfoHvALW+EkMRO/lP9fF8u4O/Vfux+
f4s+aszRuC6dyS+jmBCnRfOukRniOcd52BoFJxWMdkGEXOCYZ0xrwFwcytbDC46dbTwP2/Cfzfx2
U222dbK/uLRegdyH+B6q4mO9C8S1TuuwA07EJ9PrQoOxFymYBIswz37C3rwmMekPjY6ZxWe3iYm1
FlOr/o2zOqot2uAH5goHnFhds0BQ1d8P6DKZ6v6+kdBk8oaITwvS80EWVmP+huSEm+bR0/cX5pyl
oiXdoxHerb8jGunVGQxsst/koHUXussBY1bRgL9ov3TXxOkX0qax5ypfQ6N4q4w79MZ03WK3hetB
bInTTUbjfvaa1gi3WDGW3CaPqg9qbN2e+FY9Hz9V+LopxTUiPRtOMGj9VJXJp4pfEECtJJmkcKiW
odj1El7yMTQu0eVN9TnRPoeRPFsnLgYjn2qHhxIOBQN4p2e/h5Q/mAc6nznNzhpAgOfTJdnUS+Mx
LzqInTeby3kB69175AfodkEy2lAIpF+6+9J6TGEu3/94i3ILlvZV1iyfeJKzbOS+oZHS5Y06vCaS
RyjGLGzBeLT3M49c7TH7yWCOKGlqr1T5jhWxuQr91mlJw5GLbzCVxK7FsnPhXrfrlI5eFRENe388
bOMvCCKrLgfGyfOCt29Dly5+H0TeDX0o7qHZON4cHi5qVQOxYZQzyRMN4J2BWTGaiE/E0Rs4fz36
P7/KbxfOQUinWsuy211P3XrYeYM6MWFXj9+pn9eaZX7WDNkl+Na38LdxYjs0kBBjMqgPzCy/d9w8
VdnDzgqF8e3EY6yvtFCGLgvxJSbh5/9afpt2MYsYHi85H+SKsdV+j5h7rb1xDLPYn/GbBj0at7gz
lrYN/ktavRU+vnXAHJgx7exSY4ztn9frg66CDkfCOgFfHmLxAAEv8kfBPKS6B2aOOtyjy7dpvkL5
HplrznnAPvTJzwoxw2ZuB+SWtYSDqf+nggPnTwnJxksIuQzWhoX+uuNMSmSdnibRxgyZ3LWL6jAR
kR29CU+2Y9Nvpe5p5sE+R/7JViXz3ROQYtOTQCxtR1LhFkXf1y3KhVqCBr3IoCcgps3tWMXiaNjg
YO3at5+2aPXgLti0i9bQYE9bsJywyn63TNGPkR/EV9o18W3y68NLs5ON+jgj+/zB6IMVuoNzeX/V
4OSl3l6zwJjyzVR/u7KCYsPndle9dw/10J2iZ19GnhfYUoHR4qhZH/7WDMqqn1tFmS6FxWni/uYy
IXO+I2PwtTBJRNCxexNqv1VaKfzRhMLZ7wwn22eCinsZC7uN9HfB9gA72yQgvPa6nR/QFROMRByA
F60NlJXT98Dgqpl0uEjyAi8Dd0lByJZy36F7QWmQMDwCz7i+1dRqADAh9WV7P7/ydMQ8xH5duEcm
yTVV3mYMHqriK0lEJn+bVXaDcECfOetLebOfVIMVFpkCbBonwAIRvX2yCJ20CcLw6YlQTTlqabb7
R8fdMgm4wKXnCtnRwYQevLG4KRxJgcNk5LcIkpKfFSXi6E0N13PqXEilIIG6YW+tbGLjcSMKBLP6
wuNkGITOMJ3tWuTlTj8BHelfdCe4tcfh7mikENzDk9jdPyrMKFMZAojJ1Hqcdx7wt3aW7g3B6O2R
95pyDQvsSk/LSgUimd8VpWq+0OQRAdGEwpfMlKk4QdQdkbWripO7BcI/7yGvXGYCBPGHW2XXjmgK
3hDLVDE1g22f/T+sdNIvLfgOiFAF+EGeE27UMahCPIDuXCXl7TqmnRFRc9xzRh81FZPBbzT0ZW43
BWcIoeD5X9gud1clY6S+V2ZLn9mGsavJjWjcvaeDBjFTmdzCcHpjKUHviIY/EO4UwJMreuVfLtSe
fOjiB1P8uP7eQ6DNkaGaqb00AHyeZMfl5QdMrl/FS9pI3ryBnmrbeb/lKtF5U5lJCQYYzh1tFRIj
4xRi8yQycZJNn4n1qq+BGxR9V3PSie6BdziDIxU+1Wlc5sklB94CXVUAsyu6yfjkTxbLDFsMWuG+
cOUXl5VLGH4e3V3SLVwkzM6Z5nzFZYU/miz5Dz06f1J+10sAnWWMWy1E+gc5KH483h6Z9u/zKy4R
BYYrqAyMS/QAf+v6z8KIelClalSoB0r09RwHUSf68mV+ZVIHqPKfVn/cE4x1m7jf/Qn+agrggeVC
NNxSVvYFLtDq040mwoHzNsEWTGkAgcx1UXO+gh+z8Dy8Y7K54+aTaiUbuAtM/nFm8qmQh7TwtWw/
PToDxQ69Nz1CfOJ0nPKs2ePWrTM7oBcJdh33CYQ5XL6gatgce/UqRaYVzq+TQSmhRACBfFyleKxG
ED3icxRiMlUOIcu69FZO1u5KxxBaUYMSosgPwMVJdZcchDRJfJ3chAd0ak80Y/1duIJrR1O64PXj
CTlneCOw3azQhXDuH1dnsdKt6C49aG/sHPSbcKafCQ/XmuqF5swYDWdOdbBDT0aXCY3EbKkpWry4
iK2lEwD8RxNAOXhde9x3HnsiAPMVjn74+0H57WX5i+rDwptAI1KWe3AljDvEOHzBQ/rPmnHFO4Vr
tGT0Q8fgZKhPzUeXoEokQhbQC4GPvJidaFFgsx2b4O0O6o8SMSa4oVAcibUGXz2hYG1jZ5gZjfA2
O/LdsDUn8Ez6BpQsc4RxHJCJg82M/9Fu/MDrD/GdWFkh0FUT0isCXemH/XxrItRJn/W/h1Z65jxL
HToGeh+dyGJZ9Q0sXE3ovsIqC/8Cp6JDqVUZhW2iNe7POKbpXKNhcFn5PU+yI652pOZC5NO29nwg
NDFxT+TU5qDsvJOgsNf8QRv+Hnrp4PgQw/GPHUJE/FFYpSCXuB9IiC++oCX3bIanq1Mra+Q4MYgQ
+NXVyKk70/b/2tr5Drg5ZYkGcgjZRT8mzcRCQ698NNip0r4McAxFvBfxorKrI1Z2/4EWnLUhMoaN
nr2uYsM9XNgDJPSvqaVtwiZLJcdlpFcWA7zL5z6gO9qf53Oz+Qhiapz8sb8u28YeXVh3VJ8Vqx09
Qe+vCmBON6daM3NzVdqxWmiH1pv/tgaI+jWZQmu87HLg8sU+9Kj/CzMtdEKGAHW+dj96HD790rpU
uMvf9EyFEU7w1CtYPfEz75R4SyZdgYIY16v6Um8liWBse/xII4v72vKo1eC7cQqim6GRn4X5WRYM
FCsEOXpGIHUjVeDIKNs7QDtTxNv2j6V1jq67bEeBIeMXrYFEs/NtHMt8QUJ059yoovGEMasfMOwl
qgZ/8frW5+j9EkCbZb3tTv0qwS7l+wkV1vdiER+MUCZkq6/SvtEN+EqEVRpv/sUDnRFgWD3yzVfw
O1twR7PggfXFDwS0YS5jCTSfSq5aWmVlsbAL9bN7+Xand/yE3rJCiwP/2z9fmj/tmqhXjXpr3/ip
EzCL3NS6N2sIYbaIhPcFxZglM60G7AysJOFdVu8PKnBH7CPRUKMcKOjL1FXMM59GVzeCi9E6RGd2
5ddBjp7IhBQEKzYHkm33AHCrRX3L2h6yQ8ZV/zkSVMxZa0g35YLQjbDhixKdv7IJP1uurwPvYCMF
bwT4vks9glytGxFl4XLCjc6TS6azZ6dE+HC2zwynOqCJPjXTkejnFkuPNKZ2tFZHqOPRBn0CcqG6
oVUwLv+gOlXMsfMm0aDbJwX47aXk49l1YN2w5Z07FW84whQoGNC4+rzZchRw8Erf9lFiKtD2CPmS
pnisDaxuuP6rXSsxRzdhV1ys+hWC22402hsO/E8j6y7RT5rX7xAk4TvxYdnG/NtxhsB31JWUt+uB
+R9zuLldZeDFxyJxAMOI6USk50+kqk7IzW6/GxJlh2REsnrvZskdYQgInEHzSRqXre4kqv8ZKn8i
x6ZbCMMzrZIvaSkGBqnIvSlnm3WHtSSf+puTAbG0+VRyYdHbkGMJVt71txZIyJoUjSpmSNa9Ve9O
JFPILkIsV6kai7HNVBv2Yo6dCXFGtv9a3C7BKxnpeenUTu9FK9tabTML24hWRJpwtdmoCtHEGLOS
ouaVjK4KzOMOltboObN+JUYppwDIEguJdxgXWzTrzh7QHujJRrr+m01bY4HJ6EDPX0D3y7EHNDtB
rkR4xINSuL5YI+a4XMrevf22x7/6IGMZ1cucvJ8nwbcGK+1GBN8BeyMiUaFkjYECqCdN3iGZ7YK1
QqHGPaO/9epud764O6aWUCSUw6rw/zuGDYNyxaNMWFYBp8NVAmNLjfvlsE2021xfgYcnOAt0NQk3
3uP+mL6QKzsfsuOJDXzJ+sT9K87Mw3X1jfp+JAxiyQ9IDOn1ro1M9OTfR4UZod8Ov7tgpYrGW+iZ
V7T+HzxaQy49BsKcNFwlYlK8U4KTR8dd6QiJemFhYfi123nkkCtPZFddhkj4KB85dc6daeoEx4u6
EDsNWx4mUovW/XNCiGLw0C7qm7hGn7lRK0mfhwFJbKojuHKkPzXbkVfYbvls3J1y3VOg19O2cSEj
01t4WAYIo6Tj2zC7cjf7sKjLCh6W/BgnryzjeNVoT8PmOBTEmZTrbXpPwfr+44jY57uetKhjsKqb
z4DzKnO8zYQj1bctrS3kEACgRdrDRUzjh4OwKDMmpKnaBecZlq7vWtKj9MEYQSxd+OJkldagl4ag
0C3Q7B91gsvzoFgU7HbBkkAw1KRVKhBjo9gGfbIldtrE8WcVjs91rwNw/2XKxU9Sdzlh8fhkUqRt
DgLP2UyZodM8yw8s0/a+8QMPABVpjy92H7X7rIGA96A30ih8HamvMHnnGBMIcaAGe8oP7S0YC9LX
Mc52JY/fOe63ukfdoGpk6DhAsGeTMkvd4tKxj6NWw2pIOf+RwfrIQVXtYBv791yVrGiV/DtEh+DT
gO+YhFQ7JZ77v8E0qVVNiu+PxhS6adTbTWgg3QuGyAaEjn7nwAK4NHxIG+ENR1D7CCQcN6+wm9oT
fe0e1ogzQvTWDVRFsGh7OSzQ/QgfiXOcKH+MW6Xaooo75czeCU6nzGFdwRTS1IRGNl8jLd76GRKy
30WiCgH4DWZlAnB9pDnQA4SQ7nQjtW8CqY9ETTkd+BTJA6Q4HLcP9pe+/N1BYwWUGNz2Y2GJ9q+2
BqxqJ9st3yHhdvA37cUF3j3gbPI9NKOeVAR8nIXBOgOnD1uc9Ux1Tq03OvSgEEDjXPIk976joTk1
iHEDsK1cMfFrD0UGd3FBY8JT8rgf3m5GWVnPtE/oEtbb0AsyrR8vXe+XfypNCSuzil0Tb4rmbsEn
KT9xniSFvVEJ5hRwxwNYjSVdS5h+fWIiEmocZf9sHVR8C20KJ8oB+9TLvo5XuVBe/dlxnCOXBbgo
OV0QF7yAi5mlwsFsyW9ELOovojeMWrwiUmQE6fQbWMUihzDOl/Mn0S1cheo6YHbxbIpA4Meu2J9f
t14NgNnH3NgtS8CNPzJnNPuKrtMEhs+++7o0o7JQ04JOpBEOzjlgPrWFK/0TIiZScvTEvQxwiX5F
/uUbUd7Ae3FgKm+UiP2R6Gmegw3ewmaH8F/QgzYry5GEdMnys/Dh82WbsnQROch4xoWCqXW0hTaz
f4f4I/rRLafvfz6KcDFoX4Tl31dSRWu8+YJIuLtbHVRn3HKOlK6xF2oJLx+nAEsc9+J/Wvi5uUoc
AQbvm+cTxjZ88nIL1ZTgNT1yUSxOxFVU4K0JwL5+J3ShQ6drZScvcbGyAVYqBtBBnU3pUxy42U//
nSF7N5AoY1rl7OZRSSAhu20JPFAtvOl/MnI3nUF4dx0p5u5LXkbTefhr06nz2s2UjbRkS41tv6Ms
Y8DZSiNYGgfb3xYtL3ela2zN+VNRl/qgoEwvbSbci4LyTEpXr2TadJPHu0LWRq41as1TYtywQ9gx
wcp7y1i7nMikKzYG5FMG5p+zpHYzvkDpl1b+3gQQVCvCbyUfXBsHusIAj97Hn37hEFfrOBZScv5d
EbQ/ODD1za1hxUD8Ij554pufcLSKl8g7jbvMmKmlJNoL0uJgO5d4gTvbuSApZP+b8y9xeXEmbSKs
Ys1gXqwucYUqCyxWqBOcOyLfPL5kroROgtEXqR67V3r5i9mczR5JMhlW0YVvewgybacuyEREttv3
/YOpYYDwagdE2Xc/5IceR44TYUIf+jrOP81atZJsswG8AJejb0nOxXfeTcYUwL7ONrq9k+ITGIbF
DWFcAOnUN6EXcXjnX0T6zi6jDZHWVDmcKIQxDYg+saj4SM1g9eadHpQZzsIKnAelEhgjNS8F+N7r
F65ffL9ANqOAgC71dSQR6Ets8560dx8czAwGXlHnrFa/oUeY6YaLwqUVMlc0dy/gL2Rgcs8t0aYA
VPRy6EtfhWZjBwrxBWJyVwKnWbe+CM3T3pY1RSlOEhVo1sYvyykvZa1lFtTehShOFDn8bUoUx8ld
LPEIyzn2IBF3LYQk8iZ2iEBknoAQvWfGSdjHAk57oLo1f+zMqEli72QUYhxwCo0vGRsZMjAPuMAh
Kn2CPd6USJpF/URt2ABTcJvWfCj+i7wzzIvSB89/jvgaOtHsNoIxahtkg+AfI6oy3+VprYiStA32
r35i+F2ZoOChDml0sA5pC6NRe5zW9qLkWe8jffYgGP5oxk0/QsegXlani8KNt3xeqEUWZZItStB2
f7YC41ul67g0m89isYLdU5rGPso/mxCtPJXu/xPjZ1860+Q8mkKQAcm2H9v3Z4dr4cee82I/UQ1+
9QN2FWE2a5oKwcLiF4TkbD1N8TXAy92FAKtf6THQ0Lc0ZuorcdgRN4ng3105Ox9GTp2yJl8N0X8T
wpIlMpHMeXSF7JUfjOyuZ8+xWEo7NM2EZEpeVBzRmL+l905jbi2wxUfGn7AZDM73y1Aa+vqBJ8i3
hBRwvLBHwRjuX0o7gb/X4B0RiE7wkUzsAq9MpiRHkZHmAQVJ4seUs669umBxcSUS/iJY5pY1WM0Z
9ea6FrZNvZqVm/W6kWYEUnHrFt8eosqq0FRdqDsi8/LelyShptX5XETj8Q1IqWVrKM3vUN9nigMx
UEuuGuwXr7AhoXfkmQiKU3CfgV2iXa247xRdpIKR8Riu+zFBdkBwz11nRwjHdsFWxUEAUtLHLRql
h5H9Zc0pc4KD73EjVC9IxI7UpvxsBRviR63Is4y35ojwwemtu/rAflCBCOmeQbimrkPp+efWCWlC
hhvwNKdwBRxupIxSHzRMsU8UhLYhzFtl9023c/DpKdRkizEzMz5a/YlxSD3YeULqIxvdwBEKZ80P
FNz19nshvwJuUbcHNj15u3PemjwE9kmCXcBX+i9NM7HSGf+s/shYeupByawIqeT/1t9zlxn2AW7r
xpmkGt5fZkGN4tDVjXzvoH7ooJTXw6s+bmyYhcUMIrXL0IoYUfhGNad/azn3ius0AW6i6aYUb15p
qchKlf3ZgTM7rhsVEKT+T6r0tQepDh32Bb4CpLF1/+1lCBpnN3uGYcm5gAMkr2go503t2mMJZgsv
8XQdJPm7fgqfBbj7KCc5tVTsdZNzDYLYZApPRlprxAvTV9Cj/zclBTDG1fPhXCDnxExrs3P1XOtx
XfzFijNzkpQl4GoGemuj3hhFex/gj9ET8cu5FEaBXGPZoRFb38dQXO2ZRfo8CdN1TJmMZAerGS11
KTJJ10yZTEztna8KvjdjPQuMz7hk7zRNn4/zT5dRYDfbU6GYnWKvi+PBPqgp+QoCZTKV+7Ydtj/U
6hF13NXDMm03BQQJFIKSIvziJMZvqiXbU5qKHyOgzKUZlAQg4G730TfK+m4kCoQf5QNz5HQ3EXBX
DfQbgWwFTLuQk+MtoCWTLbU/IcYMnRxt2w+I6guk+HbaKMZ8heQ7VA5TM39w7dOYMsImwFOhQ0dw
SHrhNu841R+vU5GdNha+9K/yGxyc/X9G6E56OvhEfkFQ/eJw+w3SfuDo+y16KJKVs5RhZ6NUM1Yf
8BwqnFsZ4Pje+Pc0vSq9jcTLjyifEu9T6AajFGqi56+qt7QvlzlVelwNPlwysd0TWJKR5KLX4mrG
r2Jq4+Q6Jw+6msMRHJbEeSvYjPryYu9T+TmhtTzr6XfhB3lV7iyCZhePHgwqGMzCe+KO3AE60zrM
QTvrpZ7zUnFioYxt6t+ydx6Cy7hy29Rc2K1vny0YAkxi4UfOzd6exBXiv9QDQ6XmxZUN1A2a2wDd
3E74pcEeQVIPxOGOObKoYeT4BfA43qtkF3LZbYPbdYFPypL8T8BW6qnwM4fbS6rrLB0rorsP2Nks
jssS36pqJH8/XkTSRw6N7fpP10xPNGxk3tvW8OED2G7WkAPjDuywaOGE8Ufm2R6obScCbuVi1FRG
qLgNwt4aXVfy1ksGWcgKHiXhtoqM1M+vGKbu+I/LQ5qnofbS3twuJ1g9d4QI8ZF46jaIC7NDgAC9
eQ30/zJM5LAr5XNmP3Oronxb09Kk6wa9+YYgL8HZA90BQiXp56tqGlFBV9pDZuOjkwVVN3p5K2m7
Lu1TmMyCLquwjDuOqlPAHfyckKSLj1zqDIc7P0bOeFAzGHA+2DcLVhGh8olsf7JUG+2+xEK/STOw
WLIOJuiklG8md2UQf2Ld1kdrElGQHdWTrKm61IA8LWUAiK2NVjweSEkmfsf5wwLY9OT5w68p0qWO
UN7HlKLx50LfYrN9taVzhmobT7UInuFVreSJmJ1RQd14ihAFcdU0Xw3j9f1wy9pJSWa5Ai4TiiV9
daoz+YXBPdxlg+Ah//+ByU02QPjfN9W/jkB7ms6BnR4DcBt6lxZ7o7W5+3xcihEgDMcWIPMrnjoO
19YuIr4SgqN4DFTw0n8ym99gehwWLkH7G0V8AlknLCd52tLWwP734XHzUnFbOvzf9CSs5po+BDXZ
GRqO9LXHB5o9gJh2nUKBZe/BpIzzHDA271il40l+jnQyRJSi3NvMEEFiI9i9kM39YWsJpjqeRXJ3
Lv58VIDAItGRp9+Rm1+ITiveO6HVJ7XuT48zSga1wkzNu3JDC/0rlmdy39EzRc40oWff3NCPEwrt
q2mbKFO16/pBSRtqvLRr0DfEUSlx6TCRx5KHFhNVjhxV+oYz+f8PPQq3qzxCh8ZUR3XqplaTQkJK
CnShgCEa8aGhy71v4mrtA3gaeBEQSNGejgfBsaPfWdl0ShluTNwBph/Ne/CJtWBMMfmYISCie77c
rpTqigm1pq9mAdVS1ddofnv2pv0NEUA+s1KwdEmtipasls6++McyIAGIysskFA4FDOPJWzcjPNq6
c7kl9DYKcJZEtTzlZxa8uLOFs98QCpjxB3roIUNymF4D1mQTqYY20fkWWzgKf+b11RIUBm28LGr8
TiGUf0k/uNmsg0edp0tb1FzKS3Lrp/p3Y94nQdXJWqjiwESogWF+orjIrT6ppl8JvXjt5eICEO4X
xPoYRlss4WzQxzcHAX6fv4oB2/PTlTKGu1jbDsYTTKVMqhaARkSC04zIPkE2bbAowdoFTLjAb34Z
OAjTgQQL0O49THRHS5Ts0dg4z/rHRhSG0TxAmeKuH156biH15DTHbVVVx4yIjRqyChQWZHPANfUf
w/w5EmHZTlpveLrkyfDt84s0I9M6mQJSV50Wkwf2gOjnOmL+OtWnHT+m8wFTB7IbPmJJkAUpKHqb
DCUVmAqnHxxDBntkLWhz4SMExaTq9cUH/pYY2Wu8vtezQJz5bU7HzkqRSafqvMldEpukjgDUTHNm
xWRS4DjaJy2uA7crcIUTJc4iaN3dJ1gO48RdIuXL1ei3+Mw7s+QHyghhvxJkRYcfGlOyVRaKUmuG
0FAM+ZaOUGo8sp2i31NG1ayFvqUhAikGjcnAKk0cSximB/KOHK0JEkgxg7bC6Lx2TxX21IQG01lS
7wBrillvKklveuALDCaqt2m6BOmjJOw7uucgDBjgvFEQq8N5f6Zw53azB8WyYSLGhWzXs57K8l74
BtB1lcQ60dPcbqAraTeWrA1TpHuQgGil+qbw7VuoAETraSIq/AjZp7ZbX6eE39u3ANp5u3WhALvL
SFif4pUU1oPB4Tl+kUy4+qGp8i4wmTPyME6brdQQfIyPBSGKOFiJqT+b6RPvlr3qY16lprmizpAc
if1+edvdiY+USFZQ5mfKLgjLVcCS+DwNcxwOiOAxqIvlXEk9d2dFBhvd4ImtMgDRXJeu4rCK9BpV
Kpk9sa/sno9WcxI3xRh0cSRSvaXfqVNuoclqEv8yHdGyCg/o0nv+YspbLVnI7ueLHiuJYFTcgPXS
9+19DFMMSNVB2x+sIXqTVjpm8GdH13xRESjpBWwDJJhMZ4FdomgG1iJjHXIu7zV2EWD4Xsu7Dyfy
rMVCUnVpVJelUyWf8LoCzwUZLivVDkEp+cgXGjKDTxBPwWv6Jh88dIKaLtdDHm8pv4URGNgWntx2
ECQJoiyCoilsg+4j1wHDPVFQDjKXggHTuvQemXws/sFyJGfPng4g/t2VYlszuZiW4F0l+f4BjYKN
OFLpvbhxWXl8Mg6gfMD6KFFwQTj44UjVGOC9QJMV3pMUw9J9eDwxFrOU63pkFml4jcSt7cHo5if8
6ggQV6ds0ZjRA/svDBsYZXIuVsOLYziYHMg57nKOXxuIUZ91+j57Dv+vAIc2iLXy3eS5oyyOQons
rajgbkZmoqZttq2rIJAbSQVkqZRzmRBWeia6Ew9Yr5+NuzCYLCD+jgm0/wfTs241/QBpfBjaLcsj
WDPFSeInRt1ZG6w7JxuPE1v6MxLFVNUgM8Mk6bAqjWZD1YVTLFffOi9ILZAeBUFYURy2kjHiWs1C
xocoPHdKnv2JXfN0RnQnOyih3i062ZyK1SYn7eDNikadXFvY1Tb9XP4H5iPaNVCRYZP+vpliTIJA
v1FqhIP+U6oeEVbyZZVUcmR16SLvYuohvjQLN7Ap4/kU2bIeQnsL0PS4qMD9KZfw9wkVoUgn4FAX
lFAz8uabscJfM7elDST6u6bIK1Maca9VAbfXYUE/ylhyOvvqp/G4AKWK7/nW2CVLniobubMAkDE7
v4FLYHfYUenH4HcEoy1lArZrhpSih5G+FqjuO1/1jALje4dCzdlP2y8fEcrDQYpUnQBSpfDU+vJj
lclpgMnIllltkHuhB7A/eKosBpqzo/LwI7SwZixlYkCrhzCxRhOgNOJhcyfaIiRVQfmIc3zt0WRx
1rAD+qBUWGjNBcIsJZL7W/3V0ywpyQRMxndQqJ4CeDWtFl1B3TX8p750xIKRMEXXL0iQ0M5KNBNm
9Xrn8Avuoh6MYcusYfx3miLUCWMfpvSmhgTaCRl209glKTowRDmyB7IxFekSAwrgViuELtHWzBzO
RpqZe1mvrZpNmJJuUIZnMOtRm6v2g5cNcEoxRURENb7wmDxjYN+KDPgvH9PcwEJQp7NSnEnJ/I3p
Ii48sZIAaJK+hLBno9V6CcBPjTVYIF8Et3kesS4ob6lOS+cQ0CLKHYmwf/4NxslAnOYfEPyWFQwO
6Q2DAGTKKxHb5RRceevjWu5HPLaNcecqULahrL5SWqQdendlnp1PJLrPi6BG2sdViKeV8viVGKBE
vYYZ5tLj/tA4W91o2nSNkIwbojKmbN+AoSOwJ2M3v9tjNRfi9+aLmjOrp01J5xzZQkZy2UNYgXYo
ppgbeB633j3dHrkXx0UgqBAmWODCR1GjkFx2HXSoJ9jTvK/S3NbVm4p0cjOpDi5uo3bL1qBeomQv
gxfKiv2jOKMFLlhBWJqtcQF7qJJuGLIP2kdfIapPvck9Do85GLnNRF90b2ovBxKHtqsYl3TXdP/b
A5o2U+H54AJQF9CYh3zO4rFRESbE0ERkc/mZqmzHXOD3fWUl+g1SHndI06nrHb8N6V5pBdhhiOyX
E/IP+/jpIqWtfImd1sB6C0Zb6OGSyL8Vk7qhkjXEbLISWkcGbRsb03IM8CW3xtAWkYzVj6w6ercs
wzOg7emeVCzPjEW2KXvlSxxFAOjZsCu0imviA3bCrdD8XLDk73oIXrbnjKSgV1pWQ+6UxeUhpJcL
pKtBvFUoBe1YNHWuL3F6EExJ0bqFLGxgllf/B8H/tyK8e04GWi051u7NFtHDwJgQj1QWrChSubyW
i2cJsW6nv1zFBHMYI4Cz6ALIsbIjdc3chRp7jMeREiYoV5eSKWUcEMGsmmkGnnH8l1l+wgcML+di
pviw1rPu3Ya5ou9z+c7q+OEx4duXZDdyj/vIuvJoPblPw8pBkJP8doyITN7n5guSRw/VgZ5FhR6Y
rvBK23LDK1YUNdNY22+t7oMhGzTZYmPIKYNzNrWeMCJsxRjrq48hM5XHyBdYILPU5evwS1Wtu4r3
Q21BmALhjaarIdhU1IL/S6pTa8S93xthQv88dfqsXI6r/4Pq52boOWl1/K+eyeDuIyzmqeCzEVXo
IxOX3NjtQDA58ZK2BFvyFTCTfYuV8gK8hOXWWxPCww7BFjg9szlNeYiHmiCDtU542XUP1TUqJ1g4
vt0A1/r45jZiKYskTg9PQs5baKMjNOeX4tDLIqtLWWBZSQaHjThzqXZlALdusTf58ZA4jzuHxLwK
B+u0y+eYqdxl/1DiV+JbLuMUqmTXBQ/ltwV6Sv99HWslMIbC4M3RAatpcgdjQ3yJO7hy/BESM8FW
XTiQbDz6uBmOJTOju61XHZBWkmqyG+VbhlzhpEEGpFK6/BxrcP9r62Wjo0rUvzTzNL7GCAaews1c
1+Z2bgiF33Wd7l2JnSyvJam2F++czD64lwPkSkfhKw8ZEM8J/d7bm4m2HBD4lw288bcF+zYW6yEH
RPP3Wh3SWjjCc+mGw+eY9MJNq9sIxiyCmwpeG40cFinnbKywmphFPjk1wTzF6nFpbS8Fiu19q2p/
HIqKrXvNQvwY2YiZbl5y5y5AeU9MmAWnNUHx/tb3lXSaAoaMVx/JR2qNc+9K8KvM/Km18V3vJS/I
qzKKEQQ96fhJTuMiRQywaWcT0PKSdxiJN5QWc324ZzoIY6JiEnT2WsCHIiLVoqtOpRbP0pvcU+Q/
TpjrPd6B8eiIZQSZTwV/9lmrE+w1cnbdc2PwnQDZIJzMlTt5Ar6fh5j2Fgbu5AOnl9E/AWPPwoqY
JAsij5exGniLAx60seMsp7z+FcLSdjlIJjTS0MhV6FNKqEkNTi7ZOm4RLBQYl1/y4BkoxlHcltP6
Ju27VaFo95cc1eURbj0PSRtWafAcW5XWBdx5paHFPQD6mcPq+gPKIU1tkAJ7zqtlB3PT4MH5l/qC
UDOiIubmlEKEssLIpmrIZuXgGhPxQzrFMXSlTSsmj0frVU9c3i5gkjYfO82EKZLmH+uPwE6tPnz6
E1ps3f9824OqfCAsDgEsu/YH5lqAAj3hfljzP7TnsbhI2aBeVXIPvzQovy9HABaieOPeBX5QwwjX
bFA43Mudb+naHADgg1+4/tyXMic1G46UTsVZjIg/DO0uisRAS87FQEQPfGdvmBS0cNIjlVswDQSp
cqROARuwiX+HkOR15Py8nLp9WfsBgu269gQPoY+k6VuNucfRa82XztAAkuVgF2IG1ihayQN2utT1
R1tqX26KS/9YmO54qq+zbv+CnxzwI8B9llgZDPVzjBlXb+fclAELF2qcNh2X5PkvrtHTigOXBYmG
sT6yaJsi95uibDmoYqHDgiq+NtT8JnwkpLGQcwc4An2QfYnXs4UCfie4YAYHGLWezgColJxnNmOk
g4GtO8KDK4w2JJeFEG3FGiO8Ec8CKvsckAnArRYhjTrgn5/b7Tx174utbTpkZkfytFYW8faiGOtt
Ir0ep0zOCU3FIMf3rNoJFg0oXqBW5fuRsKFyt3wWcwFi35NZHL6GZmv7p+ue4nw5mIU/fgd+krZl
yVC90YBuen6pb/jaCAxqyGnwxPbz+A1nqIYA/k/Jlx8guEPe9uLuo9TsfqsC1Y8kXpaiIZG/2XaE
3OfjA8nXngtIw4YKHDCJ0UlfYwzyfvWqBFWJrZdmsC1ZRgV9ceUnYLMKZAvV64gO0MjZ8/i0as/e
HWQCob4gDYyPPqIfBX81cZuObV8fBbmw+K5vsQHaH+pxLe7mFtcXvzPL3cxpbcf+UZqCdjeUl57o
GRtZDv+JIvU0mbKAWYsKqLR3sv3N/uotXUkfhWLy8cqiLBenqO6DZH0ZQ26cWVarmE4xwVOQux8G
csg0W1RfsvEtpCWxEMCq3QlKTQYqLhH3lgOOJy+2/hEzM1ujNAp63KXgBGUit8lwPqtd1ecW9Bdt
lwVPRRWzoTDhZ4RzI8GpuXqmyC3bHjPJRsncoHIvMi5m2tC1ESLo83wFCKmtXmUrExBdOODzbQPs
ABQGYVhHCV7RAkdfOthh/1icl+ovaP6VdC3I9EXtq9JGqngvh4wBOtihAuXiPKeoAWfvYPCeEUeG
xseB5nLLksNlDw/QMQXt2FpSfo78vgYUrfJCkKNmMF3Sqh7ocB/4gEll26xITf2HKjevRKKNW4x2
XrZdV3bKDbmb9fBh8IIgXpHe5ZhAaBak9XotgyxQa3d/56Sir1wRXvXuasSyegDwBmldNdPGdJez
+oB5tJv1PrjEJU5WK6gkIUXKpX90J5KZr3rYp8hRK0lwlz1HNLW2/swL3TYfqw6OM1EmGczE5aTP
NkjXaIt2Svifpl2nq+QnAMfMcw86viUXA1qZznYUcXLdHLEi2yWy5Ce25RGKbbHh5A7717eJlD73
wAp+8t7FMUb9eHLr7ED8mJAYHM78Nu6/mAzAocXbdKlxD4QAE3xCUptFlfBFKr7SZ5dzFTIB6Df0
u91xEGDhccQrhosrLtuudTxnrLHxLnIG3zFcYLu5wGTs/ZO8AFnp5u1sI0BNrTuKfYyLtFCz2na1
OUh6eWosahiiUQj0V5++06sRbOLFHaENVqMGzDO0Vrig0/6Dv64Dkaxmu99ToOFyKqmYhEDcyPkh
Lcp7Al/OpTxvkeauDg5u8h2V9MD/j7d6eqxPyMDkhWCAdAdQJ1fegv5nSPaYHE5x5NZIX5St5552
Z1NnRDiJqG5kbdkFFUozHxpu288z45wXdr4xWMf6P5hDA7Qf9Vw8Q6gFQ5Ap89xEs/D+47ish3AH
oHCgN0iwbyHpfKrKi7xr/mstnwoy2rYd4BvSGj+v0lmgzg2mh25UyjXzpsNuN9RTzFVkHHC1J/IG
QuEtQpa+1JGM1eRIdFX9YkfScZFBQDI4Z/w30WL4jbMCLBGP4nRjfvI1NbtCRTvctP3WLJacy5G0
faZEG6ty7C3lK/3Nt6fSDqzAWn3oNQfVnY1Vc2cW7DI3QOWstlYWmB42UZVXcOikugeSnMTRf2SY
J/yc8U/gLq9nDvzgFluqYPfKDDlKkQOQnKss5DIGp0jysD1o23JiADRCoGTf7Y91+8izzizubOEI
283Kg62n6p8yAxWRlInf3EwhK09iAEIi8D4QqcUhxk3yOK1ExtMeUembW2u3GNgMCwxaBLpiZc64
eyEkFthi6HX7UrgZpzGFc2RaW8Zg9IlFQC95tI4V7qWpVVZ1p7T0pveOkvft3Z5mC4budyZH8CFe
uYMepemiwFmQEtcC4yEe3lwg8fIF0wSEsI9IE68ygDr++duOvj9dvmX4ZkAqVJE+ACLqQpGSUkar
BaTaC7ceBQOs2JTXabNx1no1oyxpDEVLcC6Zpn46q5SqYq9oichJOHWwG/lTxNqbk0peV9/gnqYi
408ubJmL1vhgqYVJncPEpZr8BlxO1qdBGUOpMSjLEL5tFglCXlrhl+WxeKTbm8pZyW0bGcVsUsIs
1jFreu30WJEZU6iahtBeKXmVaLl4uj21+z9jFkxZrFwHNmzKoypVIH1sztjpzRNGyux8REG1zJ9f
y4eZ8Gtks4XMOx3J9z9gyHb8K/+pFMa+p0cXVnrzes5WhmiRrmcEK2sNxgtikfnL36GlrJgPTN3s
hCjQ9Ct6WZX2ga2v0sDamsjgYisNvFI7IU9NWO2Gvj1yEA5berV75npK7tLAQTssHAClbsQQB7ge
kLk4FMSRQrM2wjCiGe0l0BfRCAV3Y08e2yLahgRqN4ahJkm9swGXgL0vg07C+JnsZkCXsLN6hkZz
3ldwIsu5Wq2EHbbqy0gzatEqwb6KtfRb4eWbmZIcNm83u+AnIzBVB5hwXHVcmh802tygIGBX6bgP
QeC8y/Qo2oflPhuOFB0dawOd1iimOcHsEqzaWxVt7MU+S64itW5PkmmxPvfmUxneKcD6M4rXXS7/
LAUSHMJNdYkZSJm+/UkYAC/GzRgKSet9jvSznZ9MqxXkpALUm8FuwOiJIf8YDy33ybHTMGbU0/CY
Zbe3WzGn0P6MP735pgzE0CtE6yfBnId6QPydf1uoWcBIU4dbe5xW6WICC49Hp/Cul0lGCV1fOQSV
s2NbGChmj+slS9OD1Daca3XD6JpdtIwxNfKSCHAm7BRlNw/fg5YlVc8QubW09LkiD+vM0wuEc0Lm
jbFhXZTXiAM2ZIIyaoqRfWYLQOIZ6Dnav1dIwqOHsVRycmOLPsiEaAND6yfIHGsARBl10gnUatSI
JVS0/hFsQKliuWP3/L7qv+By8gGQ5n2nJXoTxQGcMhxg+InhdW5uRF8QsnZPtn4QJPH+2ZvdYvfK
jndfrloqqMWAQNiYwcpDZuoKKwmHdTIvSiRNbZFY6gmh10IuKcggxMftgReBwZ/BMlCAHGVBJ6ed
MC99+WXJqH4gKPLjINAQ0WYO3rH/VwBK37Bo8P6571qiJDLstGt0isWRL8vluSI+Fqt0VO9tV1E9
v3F0B48z6/MGYxNQaqwT9R+GyL+RaAIFPOHJWTsGx70XjmroUZirbFbUpXoblQDNU0+hekI7OlPW
xS/Us6ekMByrspKw5N53tdP+NO+BN6rPi0RjzbNAwohj1NLcTESA0Ra7k6IQt+WdhR843x2vlgOl
ooYbu7C7CY/Rc2HiWRZFOTZzf+74X1/09zOTL4dq6DQZpXohvj40tIsEmwBt64zhZBLN3qXtXGBI
HjG1jPDouPplJWiFGX+Dt40cdGyUOpq4qhOdB1lcbES4YFAOZvtgSjQAtfJTtKvCADXb3wCnMDkG
F1+3Lbw4hURFUT7eSjHHjLuDaJF8V/u8fEuyuE+/Dm3J91Oxz4GZ5sHXtcHIA/fgg57ImvGJIE2T
8qwPNsAdqkAE3IuoP9H8pBUkxFMXY8AGL+O7e0yPeX7TLBM+y7OocusvxOzL1rXMrNOJq7wA312D
1iMUsh8wVLTHiwAsgby1IHTvKQ4ltFLWEq/z6ur1klfgJPjWaC7J1VBtxBeVUItB3KZyy4MgyYn8
2zn665gU9pgQRvBKtlm98hQ8kSm7UdJMu6tJe0UIyg+UiOSy7V8p355CjNb9i/CiPIbSoxi4n+XM
XaBlnMe88+5CqfYMVKSiIQ7iUug95MZtqKoyi1yNaVKVca8n1vTuhHFcxQn7xUmt/0YkWgT+zOQg
sE6o9OxirMRMWHkDoN1VX9r3S3NFPp8UR4g/w8Yuh0is/s3qKWz6gAeAgj41S+6LCmJKigovgIT3
OU6RMMgUwPp3eaZw1WuSGNa+kEunjO8YuOnWbMJpUFas52M7QABByxqU1/LnvwWy0XHIxYgIIQ9C
SB3UkS02S/EK4z0D2+3IZ+l9hzd0FV3jsYYN/7WtkJ50lNSVCvOdH7la0UruBhl6f6tq3QYN2rkE
jKrXvUSE3XJj7WmllnX/nRTve0wspOzTHB4Tkbcn1B6GE8oKcj0g/LjyiaHACyPSdoV2y5ef1Rf0
1hr7iQe1rlgxWLO+Qj8wqh6ZtWatuNBvo6BmjYE2njctJe3cLKAK7nY/67S1YT/HndWqNEY4Qgo9
mA/KgigH1E9L6U6JoUjFsg7m9nNi4yhuKOfBlxzgs2vQmvz+FYp18fquHKDLUIwJPqKP1cLpQZUB
TrBP2fXCw3duUSbthATF5ylPtN9d6u8C3SPMLpQC7UCpDxtftMvQDfBZ6A8MyHsfXoVp9s4NYAta
N4niMIqSxKUk2Z+KSEeZz1ao+Vy++jSf/uWVgInysd4XCbX8gg+bBTwo8SIbKw0tbB63ClVrGrMb
HMCfvHcsPERC6JgL2TsfdUAPjtI/H5xkXod8WjzKp7ccS6vris9cdh58gcs0CPxmsuULGD0K+V+q
TQltDe/02r34ThL7TPUAoGP3AGTvlY+XtwZmlyU2nTHJGLebXNCvn0zxiQqYPEfZwRhxq0uy6FKp
Ez5bTqIyyBPSipEdf86OBf8EW20NwBMLMTNiykHZspIlImCb8KCHbk5y/O34qMh0/30jq16okPz4
ra9WxX8UKOvCb/mbjXQ7H3itka2T3h8mSfGv+nYsR4iqyEz/0DNQC3tp62J8/cpRaWOzDbUYKN4i
wMBkJ32prftgLPkKxqClMWq6vp+Wv4B0F8wN1LwBRQUeZRNA9eDKqH9wgwcsaTlUeeH8YfxqwCsg
n71yT00cO457S51/3CgK3epXFgrubm3FuNqB8KCYfUc81ii6Rs3pjyV2La4MZVMSkqqmrl8FbPy5
tBGy6dKZEYxza19dIZTFZ1lCHwGE/qyJJXjOxLivjU5zSh0PMeZgXTKcHn1YdYactc5aLouI72zp
r3mv10LbIFfZBqt6n6PO817hu6DCNsl3JPFgrUrlYjptfngHLNl9a51STHqh2iQIgn3AeRExaexo
/cMC4woY0kUaIv1SD7sSK5L9xKXV8a02FXwDf8ieAbIX1QxOGbQoO1YvdJ/mVHUajiBP3umAbyU8
uVuU9AD8AZcRxb5zK9qPehdPWGCQmDUbcaja5ZygDtni7QG4OJ8sgJn/vBeriqzGl3qqjqtaK7QY
YMa5+ThDQ/NbktOJG++qGMvVIxNArmCxprh+blexQgLJov7WhIZ23ZlzhUbmBhpEEhmhWUSbPciq
KL0l1l7YAzdLZ6eBn+77tXuxnwG6rgzF/2+gCWuOHWvFs4p2T8PkYTzK0tfsNMPh9Q+N1Th13sw6
t1okL+ha9ltONuqoW8mfLClx4QcOAYRUt1w0ntpSZG6AE4latfiYvtZQ07rNL80zhsos6hrErXvU
a5u+Y3I2Vs8BqXGnaMWPbpoZauMbm8Y1l8BGwzNBEsa0P6wxvMAR2zOIBcxfYTVM8yhK8xpgHNd/
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity dual_video_fifo is
port(
  Data :  in std_logic_vector(31 downto 0);
  WrReset :  in std_logic;
  RdReset :  in std_logic;
  WrClk :  in std_logic;
  RdClk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  AlmostEmptyTh :  in std_logic_vector(4 downto 0);
  Almost_Empty :  out std_logic;
  Q :  out std_logic_vector(31 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end dual_video_fifo;
architecture beh of dual_video_fifo is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
component \~fifo.dual_video_fifo\
port(
  RdClk: in std_logic;
  RdReset: in std_logic;
  WrClk: in std_logic;
  WrReset: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  AlmostEmptyTh : in std_logic_vector(4 downto 0);
  Data : in std_logic_vector(31 downto 0);
  Empty: out std_logic;
  Almost_Empty: out std_logic;
  Full: out std_logic;
  Q : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_inst: \~fifo.dual_video_fifo\
port map(
  RdClk => RdClk,
  RdReset => RdReset,
  WrClk => WrClk,
  WrReset => WrReset,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  WrEn => WrEn,
  RdEn => RdEn,
  AlmostEmptyTh(4 downto 0) => AlmostEmptyTh(4 downto 0),
  Data(31 downto 0) => Data(31 downto 0),
  Empty => NN,
  Almost_Empty => Almost_Empty,
  Full => Full,
  Q(31 downto 0) => Q(31 downto 0));
  Empty <= NN;
end beh;
