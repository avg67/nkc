-- This file was generated with hex2rom written by Daniel Wallner

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gosi_rom is
	port(
		Clk	: in std_logic;
		A	: in std_logic_vector(12 downto 0);
		D	: out std_logic_vector(7 downto 0)
	);
end gosi_rom;

architecture rtl of gosi_rom is
	signal A_r : std_logic_vector(12 downto 0);
begin
	process (Clk)
	begin
		if Clk'event and Clk = '1' then
			A_r <= A;
		end if;
	end process;
	process (A_r)
	begin
		case to_integer(unsigned(A_r)) is
		when 000000 => D <= "11000011";	-- 0x0000
		when 000001 => D <= "10100011";	-- 0x0001
		when 000002 => D <= "00111111";	-- 0x0002
		when 000003 => D <= "00111010";	-- 0x0003
		when 000004 => D <= "00010110";	-- 0x0004
		when 000005 => D <= "10000000";	-- 0x0005
		when 000006 => D <= "10110111";	-- 0x0006
		when 000007 => D <= "11000000";	-- 0x0007
		when 000008 => D <= "11011011";	-- 0x0008
		when 000009 => D <= "01101000";	-- 0x0009
		when 000010 => D <= "11001011";	-- 0x000A
		when 000011 => D <= "01111111";	-- 0x000B
		when 000012 => D <= "11000010";	-- 0x000C
		when 000013 => D <= "00010101";	-- 0x000D
		when 000014 => D <= "00100000";	-- 0x000E
		when 000015 => D <= "00111110";	-- 0x000F
		when 000016 => D <= "11111111";	-- 0x0010
		when 000017 => D <= "10110111";	-- 0x0011
		when 000018 => D <= "11000011";	-- 0x0012
		when 000019 => D <= "00010110";	-- 0x0013
		when 000020 => D <= "00100000";	-- 0x0014
		when 000021 => D <= "10101111";	-- 0x0015
		when 000022 => D <= "11001001";	-- 0x0016
		when 000023 => D <= "11001101";	-- 0x0017
		when 000024 => D <= "00101001";	-- 0x0018
		when 000025 => D <= "00100000";	-- 0x0019
		when 000026 => D <= "11111110";	-- 0x001A
		when 000027 => D <= "01111011";	-- 0x001B
		when 000028 => D <= "11010010";	-- 0x001C
		when 000029 => D <= "00101000";	-- 0x001D
		when 000030 => D <= "00100000";	-- 0x001E
		when 000031 => D <= "11111110";	-- 0x001F
		when 000032 => D <= "01100001";	-- 0x0020
		when 000033 => D <= "11011010";	-- 0x0021
		when 000034 => D <= "00101000";	-- 0x0022
		when 000035 => D <= "00100000";	-- 0x0023
		when 000036 => D <= "11010110";	-- 0x0024
		when 000037 => D <= "01100001";	-- 0x0025
		when 000038 => D <= "11000110";	-- 0x0026
		when 000039 => D <= "01000001";	-- 0x0027
		when 000040 => D <= "11001001";	-- 0x0028
		when 000041 => D <= "00111010";	-- 0x0029
		when 000042 => D <= "00010110";	-- 0x002A
		when 000043 => D <= "10000000";	-- 0x002B
		when 000044 => D <= "10110111";	-- 0x002C
		when 000045 => D <= "11000010";	-- 0x002D
		when 000046 => D <= "01010001";	-- 0x002E
		when 000047 => D <= "00100000";	-- 0x002F
		when 000048 => D <= "10101111";	-- 0x0030
		when 000049 => D <= "00110010";	-- 0x0031
		when 000050 => D <= "01000101";	-- 0x0032
		when 000051 => D <= "10000000";	-- 0x0033
		when 000052 => D <= "11100101";	-- 0x0034
		when 000053 => D <= "11010101";	-- 0x0035
		when 000054 => D <= "11000101";	-- 0x0036
		when 000055 => D <= "11001101";	-- 0x0037
		when 000056 => D <= "11001100";	-- 0x0038
		when 000057 => D <= "00101100";	-- 0x0039
		when 000058 => D <= "11001101";	-- 0x003A
		when 000059 => D <= "01011001";	-- 0x003B
		when 000060 => D <= "00100000";	-- 0x003C
		when 000061 => D <= "11011011";	-- 0x003D
		when 000062 => D <= "01101000";	-- 0x003E
		when 000063 => D <= "11001011";	-- 0x003F
		when 000064 => D <= "01111111";	-- 0x0040
		when 000065 => D <= "11000010";	-- 0x0041
		when 000066 => D <= "00111010";	-- 0x0042
		when 000067 => D <= "00100000";	-- 0x0043
		when 000068 => D <= "11110101";	-- 0x0044
		when 000069 => D <= "11001101";	-- 0x0045
		when 000070 => D <= "11110000";	-- 0x0046
		when 000071 => D <= "00101100";	-- 0x0047
		when 000072 => D <= "11011011";	-- 0x0048
		when 000073 => D <= "01101001";	-- 0x0049
		when 000074 => D <= "11110001";	-- 0x004A
		when 000075 => D <= "11000001";	-- 0x004B
		when 000076 => D <= "11010001";	-- 0x004C
		when 000077 => D <= "11100001";	-- 0x004D
		when 000078 => D <= "11000011";	-- 0x004E
		when 000079 => D <= "01011000";	-- 0x004F
		when 000080 => D <= "00100000";	-- 0x0050
		when 000081 => D <= "10101111";	-- 0x0051
		when 000082 => D <= "00110010";	-- 0x0052
		when 000083 => D <= "00010110";	-- 0x0053
		when 000084 => D <= "10000000";	-- 0x0054
		when 000085 => D <= "00111010";	-- 0x0055
		when 000086 => D <= "00010111";	-- 0x0056
		when 000087 => D <= "10000000";	-- 0x0057
		when 000088 => D <= "11001001";	-- 0x0058
		when 000089 => D <= "00111010";	-- 0x0059
		when 000090 => D <= "00100101";	-- 0x005A
		when 000091 => D <= "10000000";	-- 0x005B
		when 000092 => D <= "10110111";	-- 0x005C
		when 000093 => D <= "11001010";	-- 0x005D
		when 000094 => D <= "10001010";	-- 0x005E
		when 000095 => D <= "00100000";	-- 0x005F
		when 000096 => D <= "11001101";	-- 0x0060
		when 000097 => D <= "01010000";	-- 0x0061
		when 000098 => D <= "00100010";	-- 0x0062
		when 000099 => D <= "11011010";	-- 0x0063
		when 000100 => D <= "10001010";	-- 0x0064
		when 000101 => D <= "00100000";	-- 0x0065
		when 000102 => D <= "11001101";	-- 0x0066
		when 000103 => D <= "00011001";	-- 0x0067
		when 000104 => D <= "00100101";	-- 0x0068
		when 000105 => D <= "00111010";	-- 0x0069
		when 000106 => D <= "00100110";	-- 0x006A
		when 000107 => D <= "10000000";	-- 0x006B
		when 000108 => D <= "11111110";	-- 0x006C
		when 000109 => D <= "00000001";	-- 0x006D
		when 000110 => D <= "11000010";	-- 0x006E
		when 000111 => D <= "10000110";	-- 0x006F
		when 000112 => D <= "00100000";	-- 0x0070
		when 000113 => D <= "00111010";	-- 0x0071
		when 000114 => D <= "00100101";	-- 0x0072
		when 000115 => D <= "10000000";	-- 0x0073
		when 000116 => D <= "00110010";	-- 0x0074
		when 000117 => D <= "00100110";	-- 0x0075
		when 000118 => D <= "10000000";	-- 0x0076
		when 000119 => D <= "00111010";	-- 0x0077
		when 000120 => D <= "01000101";	-- 0x0078
		when 000121 => D <= "10000000";	-- 0x0079
		when 000122 => D <= "00111100";	-- 0x007A
		when 000123 => D <= "11100110";	-- 0x007B
		when 000124 => D <= "00000011";	-- 0x007C
		when 000125 => D <= "00110010";	-- 0x007D
		when 000126 => D <= "01000101";	-- 0x007E
		when 000127 => D <= "10000000";	-- 0x007F
		when 000128 => D <= "11001101";	-- 0x0080
		when 000129 => D <= "01011000";	-- 0x0081
		when 000130 => D <= "00100001";	-- 0x0082
		when 000131 => D <= "11000011";	-- 0x0083
		when 000132 => D <= "10001010";	-- 0x0084
		when 000133 => D <= "00100000";	-- 0x0085
		when 000134 => D <= "00111101";	-- 0x0086
		when 000135 => D <= "00110010";	-- 0x0087
		when 000136 => D <= "00100110";	-- 0x0088
		when 000137 => D <= "10000000";	-- 0x0089
		when 000138 => D <= "00111010";	-- 0x008A
		when 000139 => D <= "00100111";	-- 0x008B
		when 000140 => D <= "10000000";	-- 0x008C
		when 000141 => D <= "10110111";	-- 0x008D
		when 000142 => D <= "11001010";	-- 0x008E
		when 000143 => D <= "10111100";	-- 0x008F
		when 000144 => D <= "00100000";	-- 0x0090
		when 000145 => D <= "11001101";	-- 0x0091
		when 000146 => D <= "01010000";	-- 0x0092
		when 000147 => D <= "00100010";	-- 0x0093
		when 000148 => D <= "11011010";	-- 0x0094
		when 000149 => D <= "10111100";	-- 0x0095
		when 000150 => D <= "00100000";	-- 0x0096
		when 000151 => D <= "11001101";	-- 0x0097
		when 000152 => D <= "00011001";	-- 0x0098
		when 000153 => D <= "00100101";	-- 0x0099
		when 000154 => D <= "00111010";	-- 0x009A
		when 000155 => D <= "00101000";	-- 0x009B
		when 000156 => D <= "10000000";	-- 0x009C
		when 000157 => D <= "11111110";	-- 0x009D
		when 000158 => D <= "00000001";	-- 0x009E
		when 000159 => D <= "11000010";	-- 0x009F
		when 000160 => D <= "10111000";	-- 0x00A0
		when 000161 => D <= "00100000";	-- 0x00A1
		when 000162 => D <= "00111010";	-- 0x00A2
		when 000163 => D <= "00100111";	-- 0x00A3
		when 000164 => D <= "10000000";	-- 0x00A4
		when 000165 => D <= "00110010";	-- 0x00A5
		when 000166 => D <= "00101000";	-- 0x00A6
		when 000167 => D <= "10000000";	-- 0x00A7
		when 000168 => D <= "00111010";	-- 0x00A8
		when 000169 => D <= "01000101";	-- 0x00A9
		when 000170 => D <= "10000000";	-- 0x00AA
		when 000171 => D <= "11101110";	-- 0x00AB
		when 000172 => D <= "00000001";	-- 0x00AC
		when 000173 => D <= "11100110";	-- 0x00AD
		when 000174 => D <= "00000011";	-- 0x00AE
		when 000175 => D <= "00110010";	-- 0x00AF
		when 000176 => D <= "01000101";	-- 0x00B0
		when 000177 => D <= "10000000";	-- 0x00B1
		when 000178 => D <= "11001101";	-- 0x00B2
		when 000179 => D <= "01011000";	-- 0x00B3
		when 000180 => D <= "00100001";	-- 0x00B4
		when 000181 => D <= "11000011";	-- 0x00B5
		when 000182 => D <= "10111100";	-- 0x00B6
		when 000183 => D <= "00100000";	-- 0x00B7
		when 000184 => D <= "00111101";	-- 0x00B8
		when 000185 => D <= "00110010";	-- 0x00B9
		when 000186 => D <= "00101000";	-- 0x00BA
		when 000187 => D <= "10000000";	-- 0x00BB
		when 000188 => D <= "11001001";	-- 0x00BC
		when 000189 => D <= "00111110";	-- 0x00BD
		when 000190 => D <= "01010011";	-- 0x00BE
		when 000191 => D <= "11010011";	-- 0x00BF
		when 000192 => D <= "11001010";	-- 0x00C0
		when 000193 => D <= "00111110";	-- 0x00C1
		when 000194 => D <= "01010000";	-- 0x00C2
		when 000195 => D <= "11010011";	-- 0x00C3
		when 000196 => D <= "11001010";	-- 0x00C4
		when 000197 => D <= "11001001";	-- 0x00C5
		when 000198 => D <= "11011011";	-- 0x00C6
		when 000199 => D <= "11001010";	-- 0x00C7
		when 000200 => D <= "11100110";	-- 0x00C8
		when 000201 => D <= "00000001";	-- 0x00C9
		when 000202 => D <= "00101000";	-- 0x00CA
		when 000203 => D <= "11111010";	-- 0x00CB
		when 000204 => D <= "11011011";	-- 0x00CC
		when 000205 => D <= "11001011";	-- 0x00CD
		when 000206 => D <= "11001001";	-- 0x00CE
		when 000207 => D <= "11011011";	-- 0x00CF
		when 000208 => D <= "11001010";	-- 0x00D0
		when 000209 => D <= "11100110";	-- 0x00D1
		when 000210 => D <= "00000010";	-- 0x00D2
		when 000211 => D <= "00101000";	-- 0x00D3
		when 000212 => D <= "11111010";	-- 0x00D4
		when 000213 => D <= "01111001";	-- 0x00D5
		when 000214 => D <= "11010011";	-- 0x00D6
		when 000215 => D <= "11001011";	-- 0x00D7
		when 000216 => D <= "11001001";	-- 0x00D8
		when 000217 => D <= "11011011";	-- 0x00D9
		when 000218 => D <= "01001001";	-- 0x00DA
		when 000219 => D <= "00001111";	-- 0x00DB
		when 000220 => D <= "00111000";	-- 0x00DC
		when 000221 => D <= "11111011";	-- 0x00DD
		when 000222 => D <= "01111001";	-- 0x00DE
		when 000223 => D <= "11010011";	-- 0x00DF
		when 000224 => D <= "01001000";	-- 0x00E0
		when 000225 => D <= "10101111";	-- 0x00E1
		when 000226 => D <= "11010011";	-- 0x00E2
		when 000227 => D <= "01001001";	-- 0x00E3
		when 000228 => D <= "00111110";	-- 0x00E4
		when 000229 => D <= "00000001";	-- 0x00E5
		when 000230 => D <= "11010011";	-- 0x00E6
		when 000231 => D <= "01001001";	-- 0x00E7
		when 000232 => D <= "01111001";	-- 0x00E8
		when 000233 => D <= "11001001";	-- 0x00E9
		when 000234 => D <= "11110101";	-- 0x00EA
		when 000235 => D <= "11011011";	-- 0x00EB
		when 000236 => D <= "01110000";	-- 0x00EC
		when 000237 => D <= "11100110";	-- 0x00ED
		when 000238 => D <= "00000100";	-- 0x00EE
		when 000239 => D <= "00101000";	-- 0x00EF
		when 000240 => D <= "11111010";	-- 0x00F0
		when 000241 => D <= "11110001";	-- 0x00F1
		when 000242 => D <= "11001001";	-- 0x00F2
		when 000243 => D <= "11001101";	-- 0x00F3
		when 000244 => D <= "11101010";	-- 0x00F4
		when 000245 => D <= "00100000";	-- 0x00F5
		when 000246 => D <= "11010011";	-- 0x00F6
		when 000247 => D <= "01110000";	-- 0x00F7
		when 000248 => D <= "11001001";	-- 0x00F8
		when 000249 => D <= "11001101";	-- 0x00F9
		when 000250 => D <= "11101010";	-- 0x00FA
		when 000251 => D <= "00100000";	-- 0x00FB
		when 000252 => D <= "11100110";	-- 0x00FC
		when 000253 => D <= "11110000";	-- 0x00FD
		when 000254 => D <= "11010011";	-- 0x00FE
		when 000255 => D <= "01100000";	-- 0x00FF
		when 000256 => D <= "00111110";	-- 0x0100
		when 000257 => D <= "00000111";	-- 0x0101
		when 000258 => D <= "11010011";	-- 0x0102
		when 000259 => D <= "01110001";	-- 0x0103
		when 000260 => D <= "00111110";	-- 0x0104
		when 000261 => D <= "00000100";	-- 0x0105
		when 000262 => D <= "11001101";	-- 0x0106
		when 000263 => D <= "11110011";	-- 0x0107
		when 000264 => D <= "00100000";	-- 0x0108
		when 000265 => D <= "11001101";	-- 0x0109
		when 000266 => D <= "11101010";	-- 0x010A
		when 000267 => D <= "00100000";	-- 0x010B
		when 000268 => D <= "00111110";	-- 0x010C
		when 000269 => D <= "00000011";	-- 0x010D
		when 000270 => D <= "11010011";	-- 0x010E
		when 000271 => D <= "01110001";	-- 0x010F
		when 000272 => D <= "11001001";	-- 0x0110
		when 000273 => D <= "00111110";	-- 0x0111
		when 000274 => D <= "00000000";	-- 0x0112
		when 000275 => D <= "11001101";	-- 0x0113
		when 000276 => D <= "11111001";	-- 0x0114
		when 000277 => D <= "00100000";	-- 0x0115
		when 000278 => D <= "00111110";	-- 0x0116
		when 000279 => D <= "01010000";	-- 0x0117
		when 000280 => D <= "11001101";	-- 0x0118
		when 000281 => D <= "11111001";	-- 0x0119
		when 000282 => D <= "00100000";	-- 0x011A
		when 000283 => D <= "00111110";	-- 0x011B
		when 000284 => D <= "10100000";	-- 0x011C
		when 000285 => D <= "11001101";	-- 0x011D
		when 000286 => D <= "11111001";	-- 0x011E
		when 000287 => D <= "00100000";	-- 0x011F
		when 000288 => D <= "00111110";	-- 0x0120
		when 000289 => D <= "11110000";	-- 0x0121
		when 000290 => D <= "11001101";	-- 0x0122
		when 000291 => D <= "11111001";	-- 0x0123
		when 000292 => D <= "00100000";	-- 0x0124
		when 000293 => D <= "00100001";	-- 0x0125
		when 000294 => D <= "01011010";	-- 0x0126
		when 000295 => D <= "10000000";	-- 0x0127
		when 000296 => D <= "00010001";	-- 0x0128
		when 000297 => D <= "01011011";	-- 0x0129
		when 000298 => D <= "10000000";	-- 0x012A
		when 000299 => D <= "00000001";	-- 0x012B
		when 000300 => D <= "01111111";	-- 0x012C
		when 000301 => D <= "00000010";	-- 0x012D
		when 000302 => D <= "00110110";	-- 0x012E
		when 000303 => D <= "00100000";	-- 0x012F
		when 000304 => D <= "11101101";	-- 0x0130
		when 000305 => D <= "10110000";	-- 0x0131
		when 000306 => D <= "10101111";	-- 0x0132
		when 000307 => D <= "00110010";	-- 0x0133
		when 000308 => D <= "01001000";	-- 0x0134
		when 000309 => D <= "10000000";	-- 0x0135
		when 000310 => D <= "00110010";	-- 0x0136
		when 000311 => D <= "01001001";	-- 0x0137
		when 000312 => D <= "10000000";	-- 0x0138
		when 000313 => D <= "00100001";	-- 0x0139
		when 000314 => D <= "01010010";	-- 0x013A
		when 000315 => D <= "10000000";	-- 0x013B
		when 000316 => D <= "00001110";	-- 0x013C
		when 000317 => D <= "00000000";	-- 0x013D
		when 000318 => D <= "00000110";	-- 0x013E
		when 000319 => D <= "00001000";	-- 0x013F
		when 000320 => D <= "01110001";	-- 0x0140
		when 000321 => D <= "00001100";	-- 0x0141
		when 000322 => D <= "00100011";	-- 0x0142
		when 000323 => D <= "00000101";	-- 0x0143
		when 000324 => D <= "11000010";	-- 0x0144
		when 000325 => D <= "01000000";	-- 0x0145
		when 000326 => D <= "00100001";	-- 0x0146
		when 000327 => D <= "00100001";	-- 0x0147
		when 000328 => D <= "01001010";	-- 0x0148
		when 000329 => D <= "10000000";	-- 0x0149
		when 000330 => D <= "00000110";	-- 0x014A
		when 000331 => D <= "00001000";	-- 0x014B
		when 000332 => D <= "00110110";	-- 0x014C
		when 000333 => D <= "00000000";	-- 0x014D
		when 000334 => D <= "00100011";	-- 0x014E
		when 000335 => D <= "00000101";	-- 0x014F
		when 000336 => D <= "11000010";	-- 0x0150
		when 000337 => D <= "01001100";	-- 0x0151
		when 000338 => D <= "00100001";	-- 0x0152
		when 000339 => D <= "10101111";	-- 0x0153
		when 000340 => D <= "00110010";	-- 0x0154
		when 000341 => D <= "00101001";	-- 0x0155
		when 000342 => D <= "10000000";	-- 0x0156
		when 000343 => D <= "11001001";	-- 0x0157
		when 000344 => D <= "00111010";	-- 0x0158
		when 000345 => D <= "01000110";	-- 0x0159
		when 000346 => D <= "10000000";	-- 0x015A
		when 000347 => D <= "00000111";	-- 0x015B
		when 000348 => D <= "00000111";	-- 0x015C
		when 000349 => D <= "11100110";	-- 0x015D
		when 000350 => D <= "00001100";	-- 0x015E
		when 000351 => D <= "01000111";	-- 0x015F
		when 000352 => D <= "00111010";	-- 0x0160
		when 000353 => D <= "01000101";	-- 0x0161
		when 000354 => D <= "10000000";	-- 0x0162
		when 000355 => D <= "11100110";	-- 0x0163
		when 000356 => D <= "00000011";	-- 0x0164
		when 000357 => D <= "10110000";	-- 0x0165
		when 000358 => D <= "00000111";	-- 0x0166
		when 000359 => D <= "00000111";	-- 0x0167
		when 000360 => D <= "00000111";	-- 0x0168
		when 000361 => D <= "00000111";	-- 0x0169
		when 000362 => D <= "11001101";	-- 0x016A
		when 000363 => D <= "11101010";	-- 0x016B
		when 000364 => D <= "00100000";	-- 0x016C
		when 000365 => D <= "11000101";	-- 0x016D
		when 000366 => D <= "11100110";	-- 0x016E
		when 000367 => D <= "11110000";	-- 0x016F
		when 000368 => D <= "01000111";	-- 0x0170
		when 000369 => D <= "11011011";	-- 0x0171
		when 000370 => D <= "01100000";	-- 0x0172
		when 000371 => D <= "11100110";	-- 0x0173
		when 000372 => D <= "00001111";	-- 0x0174
		when 000373 => D <= "10110000";	-- 0x0175
		when 000374 => D <= "11010011";	-- 0x0176
		when 000375 => D <= "01100000";	-- 0x0177
		when 000376 => D <= "11000001";	-- 0x0178
		when 000377 => D <= "11001001";	-- 0x0179
		when 000378 => D <= "11001101";	-- 0x017A
		when 000379 => D <= "11101010";	-- 0x017B
		when 000380 => D <= "00100000";	-- 0x017C
		when 000381 => D <= "01111100";	-- 0x017D
		when 000382 => D <= "11010011";	-- 0x017E
		when 000383 => D <= "01111000";	-- 0x017F
		when 000384 => D <= "01111101";	-- 0x0180
		when 000385 => D <= "11010011";	-- 0x0181
		when 000386 => D <= "01111001";	-- 0x0182
		when 000387 => D <= "01111010";	-- 0x0183
		when 000388 => D <= "11010011";	-- 0x0184
		when 000389 => D <= "01111010";	-- 0x0185
		when 000390 => D <= "01111011";	-- 0x0186
		when 000391 => D <= "11010011";	-- 0x0187
		when 000392 => D <= "01111011";	-- 0x0188
		when 000393 => D <= "11001001";	-- 0x0189
		when 000394 => D <= "00100010";	-- 0x018A
		when 000395 => D <= "00011000";	-- 0x018B
		when 000396 => D <= "10000000";	-- 0x018C
		when 000397 => D <= "11101101";	-- 0x018D
		when 000398 => D <= "01010011";	-- 0x018E
		when 000399 => D <= "00011010";	-- 0x018F
		when 000400 => D <= "10000000";	-- 0x0190
		when 000401 => D <= "11001101";	-- 0x0191
		when 000402 => D <= "11101010";	-- 0x0192
		when 000403 => D <= "00100000";	-- 0x0193
		when 000404 => D <= "11011011";	-- 0x0194
		when 000405 => D <= "01111000";	-- 0x0195
		when 000406 => D <= "11001011";	-- 0x0196
		when 000407 => D <= "01011111";	-- 0x0197
		when 000408 => D <= "00101000";	-- 0x0198
		when 000409 => D <= "00000010";	-- 0x0199
		when 000410 => D <= "11110110";	-- 0x019A
		when 000411 => D <= "11110000";	-- 0x019B
		when 000412 => D <= "01010111";	-- 0x019C
		when 000413 => D <= "11011011";	-- 0x019D
		when 000414 => D <= "01111001";	-- 0x019E
		when 000415 => D <= "01011111";	-- 0x019F
		when 000416 => D <= "11101101";	-- 0x01A0
		when 000417 => D <= "01010011";	-- 0x01A1
		when 000418 => D <= "00011100";	-- 0x01A2
		when 000419 => D <= "10000000";	-- 0x01A3
		when 000420 => D <= "00101010";	-- 0x01A4
		when 000421 => D <= "00011000";	-- 0x01A5
		when 000422 => D <= "10000000";	-- 0x01A6
		when 000423 => D <= "10101111";	-- 0x01A7
		when 000424 => D <= "11101101";	-- 0x01A8
		when 000425 => D <= "01010010";	-- 0x01A9
		when 000426 => D <= "00100010";	-- 0x01AA
		when 000427 => D <= "00100000";	-- 0x01AB
		when 000428 => D <= "10000000";	-- 0x01AC
		when 000429 => D <= "11011011";	-- 0x01AD
		when 000430 => D <= "01111010";	-- 0x01AE
		when 000431 => D <= "11001011";	-- 0x01AF
		when 000432 => D <= "01011111";	-- 0x01B0
		when 000433 => D <= "00101000";	-- 0x01B1
		when 000434 => D <= "00000010";	-- 0x01B2
		when 000435 => D <= "11110110";	-- 0x01B3
		when 000436 => D <= "11110000";	-- 0x01B4
		when 000437 => D <= "01010111";	-- 0x01B5
		when 000438 => D <= "11011011";	-- 0x01B6
		when 000439 => D <= "01111011";	-- 0x01B7
		when 000440 => D <= "01011111";	-- 0x01B8
		when 000441 => D <= "11101101";	-- 0x01B9
		when 000442 => D <= "01010011";	-- 0x01BA
		when 000443 => D <= "00011110";	-- 0x01BB
		when 000444 => D <= "10000000";	-- 0x01BC
		when 000445 => D <= "00101010";	-- 0x01BD
		when 000446 => D <= "00011010";	-- 0x01BE
		when 000447 => D <= "10000000";	-- 0x01BF
		when 000448 => D <= "10101111";	-- 0x01C0
		when 000449 => D <= "11101101";	-- 0x01C1
		when 000450 => D <= "01010010";	-- 0x01C2
		when 000451 => D <= "00100010";	-- 0x01C3
		when 000452 => D <= "00100010";	-- 0x01C4
		when 000453 => D <= "10000000";	-- 0x01C5
		when 000454 => D <= "11101101";	-- 0x01C6
		when 000455 => D <= "01011011";	-- 0x01C7
		when 000456 => D <= "00100000";	-- 0x01C8
		when 000457 => D <= "10000000";	-- 0x01C9
		when 000458 => D <= "11001011";	-- 0x01CA
		when 000459 => D <= "01111100";	-- 0x01CB
		when 000460 => D <= "00101000";	-- 0x01CC
		when 000461 => D <= "00000011";	-- 0x01CD
		when 000462 => D <= "11001101";	-- 0x01CE
		when 000463 => D <= "11111010";	-- 0x01CF
		when 000464 => D <= "00100010";	-- 0x01D0
		when 000465 => D <= "11001011";	-- 0x01D1
		when 000466 => D <= "01111010";	-- 0x01D2
		when 000467 => D <= "00101000";	-- 0x01D3
		when 000468 => D <= "00000101";	-- 0x01D4
		when 000469 => D <= "11101011";	-- 0x01D5
		when 000470 => D <= "11001101";	-- 0x01D6
		when 000471 => D <= "11111010";	-- 0x01D7
		when 000472 => D <= "00100010";	-- 0x01D8
		when 000473 => D <= "11101011";	-- 0x01D9
		when 000474 => D <= "01111100";	-- 0x01DA
		when 000475 => D <= "10110111";	-- 0x01DB
		when 000476 => D <= "11000010";	-- 0x01DC
		when 000477 => D <= "11100100";	-- 0x01DD
		when 000478 => D <= "00100001";	-- 0x01DE
		when 000479 => D <= "01111010";	-- 0x01DF
		when 000480 => D <= "10110111";	-- 0x01E0
		when 000481 => D <= "11001010";	-- 0x01E1
		when 000482 => D <= "00010011";	-- 0x01E2
		when 000483 => D <= "00100010";	-- 0x01E3
		when 000484 => D <= "00101010";	-- 0x01E4
		when 000485 => D <= "00011000";	-- 0x01E5
		when 000486 => D <= "10000000";	-- 0x01E6
		when 000487 => D <= "11101101";	-- 0x01E7
		when 000488 => D <= "01011011";	-- 0x01E8
		when 000489 => D <= "00011010";	-- 0x01E9
		when 000490 => D <= "10000000";	-- 0x01EA
		when 000491 => D <= "11100101";	-- 0x01EB
		when 000492 => D <= "11010101";	-- 0x01EC
		when 000493 => D <= "00101010";	-- 0x01ED
		when 000494 => D <= "00100000";	-- 0x01EE
		when 000495 => D <= "10000000";	-- 0x01EF
		when 000496 => D <= "11001011";	-- 0x01F0
		when 000497 => D <= "00101100";	-- 0x01F1
		when 000498 => D <= "11001011";	-- 0x01F2
		when 000499 => D <= "00011101";	-- 0x01F3
		when 000500 => D <= "11101101";	-- 0x01F4
		when 000501 => D <= "01011011";	-- 0x01F5
		when 000502 => D <= "00011100";	-- 0x01F6
		when 000503 => D <= "10000000";	-- 0x01F7
		when 000504 => D <= "00011001";	-- 0x01F8
		when 000505 => D <= "11100101";	-- 0x01F9
		when 000506 => D <= "00101010";	-- 0x01FA
		when 000507 => D <= "00100010";	-- 0x01FB
		when 000508 => D <= "10000000";	-- 0x01FC
		when 000509 => D <= "11001011";	-- 0x01FD
		when 000510 => D <= "00101100";	-- 0x01FE
		when 000511 => D <= "11001011";	-- 0x01FF
		when 000512 => D <= "00011101";	-- 0x0200
		when 000513 => D <= "11101101";	-- 0x0201
		when 000514 => D <= "01011011";	-- 0x0202
		when 000515 => D <= "00011110";	-- 0x0203
		when 000516 => D <= "10000000";	-- 0x0204
		when 000517 => D <= "00011001";	-- 0x0205
		when 000518 => D <= "11101011";	-- 0x0206
		when 000519 => D <= "11100001";	-- 0x0207
		when 000520 => D <= "11001101";	-- 0x0208
		when 000521 => D <= "10001010";	-- 0x0209
		when 000522 => D <= "00100001";	-- 0x020A
		when 000523 => D <= "11010001";	-- 0x020B
		when 000524 => D <= "11100001";	-- 0x020C
		when 000525 => D <= "11001101";	-- 0x020D
		when 000526 => D <= "10001010";	-- 0x020E
		when 000527 => D <= "00100001";	-- 0x020F
		when 000528 => D <= "11000011";	-- 0x0210
		when 000529 => D <= "00011101";	-- 0x0211
		when 000530 => D <= "00100010";	-- 0x0212
		when 000531 => D <= "00101010";	-- 0x0213
		when 000532 => D <= "00100000";	-- 0x0214
		when 000533 => D <= "10000000";	-- 0x0215
		when 000534 => D <= "11101101";	-- 0x0216
		when 000535 => D <= "01011011";	-- 0x0217
		when 000536 => D <= "00100010";	-- 0x0218
		when 000537 => D <= "10000000";	-- 0x0219
		when 000538 => D <= "11001101";	-- 0x021A
		when 000539 => D <= "00011110";	-- 0x021B
		when 000540 => D <= "00100010";	-- 0x021C
		when 000541 => D <= "11001001";	-- 0x021D
		when 000542 => D <= "00000110";	-- 0x021E
		when 000543 => D <= "00010001";	-- 0x021F
		when 000544 => D <= "11001011";	-- 0x0220
		when 000545 => D <= "01111100";	-- 0x0221
		when 000546 => D <= "00101000";	-- 0x0222
		when 000547 => D <= "00000101";	-- 0x0223
		when 000548 => D <= "11001101";	-- 0x0224
		when 000549 => D <= "11111010";	-- 0x0225
		when 000550 => D <= "00100010";	-- 0x0226
		when 000551 => D <= "11001011";	-- 0x0227
		when 000552 => D <= "11001000";	-- 0x0228
		when 000553 => D <= "11001011";	-- 0x0229
		when 000554 => D <= "01111010";	-- 0x022A
		when 000555 => D <= "00101000";	-- 0x022B
		when 000556 => D <= "00000111";	-- 0x022C
		when 000557 => D <= "11101011";	-- 0x022D
		when 000558 => D <= "11001101";	-- 0x022E
		when 000559 => D <= "11111010";	-- 0x022F
		when 000560 => D <= "00100010";	-- 0x0230
		when 000561 => D <= "11101011";	-- 0x0231
		when 000562 => D <= "11001011";	-- 0x0232
		when 000563 => D <= "11010000";	-- 0x0233
		when 000564 => D <= "11001101";	-- 0x0234
		when 000565 => D <= "11101010";	-- 0x0235
		when 000566 => D <= "00100000";	-- 0x0236
		when 000567 => D <= "01111101";	-- 0x0237
		when 000568 => D <= "11010011";	-- 0x0238
		when 000569 => D <= "01110101";	-- 0x0239
		when 000570 => D <= "01111011";	-- 0x023A
		when 000571 => D <= "11010011";	-- 0x023B
		when 000572 => D <= "01110111";	-- 0x023C
		when 000573 => D <= "01111000";	-- 0x023D
		when 000574 => D <= "11001101";	-- 0x023E
		when 000575 => D <= "11110011";	-- 0x023F
		when 000576 => D <= "00100000";	-- 0x0240
		when 000577 => D <= "11001001";	-- 0x0241
		when 000578 => D <= "00111110";	-- 0x0242
		when 000579 => D <= "00000000";	-- 0x0243
		when 000580 => D <= "00011000";	-- 0x0244
		when 000581 => D <= "00000010";	-- 0x0245
		when 000582 => D <= "00111110";	-- 0x0246
		when 000583 => D <= "00000001";	-- 0x0247
		when 000584 => D <= "11001101";	-- 0x0248
		when 000585 => D <= "11110011";	-- 0x0249
		when 000586 => D <= "00100000";	-- 0x024A
		when 000587 => D <= "00111110";	-- 0x024B
		when 000588 => D <= "00000010";	-- 0x024C
		when 000589 => D <= "11000011";	-- 0x024D
		when 000590 => D <= "11110011";	-- 0x024E
		when 000591 => D <= "00100000";	-- 0x024F
		when 000592 => D <= "11011011";	-- 0x0250
		when 000593 => D <= "01110000";	-- 0x0251
		when 000594 => D <= "11100110";	-- 0x0252
		when 000595 => D <= "00000010";	-- 0x0253
		when 000596 => D <= "00101000";	-- 0x0254
		when 000597 => D <= "00001100";	-- 0x0255
		when 000598 => D <= "00111010";	-- 0x0256
		when 000599 => D <= "00101010";	-- 0x0257
		when 000600 => D <= "10000000";	-- 0x0258
		when 000601 => D <= "10110111";	-- 0x0259
		when 000602 => D <= "00110111";	-- 0x025A
		when 000603 => D <= "11000000";	-- 0x025B
		when 000604 => D <= "00111100";	-- 0x025C
		when 000605 => D <= "00110010";	-- 0x025D
		when 000606 => D <= "00101010";	-- 0x025E
		when 000607 => D <= "10000000";	-- 0x025F
		when 000608 => D <= "10101111";	-- 0x0260
		when 000609 => D <= "11001001";	-- 0x0261
		when 000610 => D <= "10101111";	-- 0x0262
		when 000611 => D <= "00110010";	-- 0x0263
		when 000612 => D <= "00101010";	-- 0x0264
		when 000613 => D <= "10000000";	-- 0x0265
		when 000614 => D <= "00110111";	-- 0x0266
		when 000615 => D <= "11001001";	-- 0x0267
		when 000616 => D <= "11001101";	-- 0x0268
		when 000617 => D <= "11101010";	-- 0x0269
		when 000618 => D <= "00100000";	-- 0x026A
		when 000619 => D <= "11010011";	-- 0x026B
		when 000620 => D <= "01110011";	-- 0x026C
		when 000621 => D <= "11001001";	-- 0x026D
		when 000622 => D <= "11001101";	-- 0x026E
		when 000623 => D <= "11101010";	-- 0x026F
		when 000624 => D <= "00100000";	-- 0x0270
		when 000625 => D <= "11010011";	-- 0x0271
		when 000626 => D <= "01110010";	-- 0x0272
		when 000627 => D <= "11001001";	-- 0x0273
		when 000628 => D <= "11001101";	-- 0x0274
		when 000629 => D <= "01000110";	-- 0x0275
		when 000630 => D <= "00100010";	-- 0x0276
		when 000631 => D <= "00111110";	-- 0x0277
		when 000632 => D <= "00000000";	-- 0x0278
		when 000633 => D <= "11001101";	-- 0x0279
		when 000634 => D <= "01101000";	-- 0x027A
		when 000635 => D <= "00100010";	-- 0x027B
		when 000636 => D <= "00111110";	-- 0x027C
		when 000637 => D <= "00000000";	-- 0x027D
		when 000638 => D <= "11001101";	-- 0x027E
		when 000639 => D <= "01101110";	-- 0x027F
		when 000640 => D <= "00100010";	-- 0x0280
		when 000641 => D <= "00010001";	-- 0x0281
		when 000642 => D <= "00000000";	-- 0x0282
		when 000643 => D <= "00000000";	-- 0x0283
		when 000644 => D <= "00000110";	-- 0x0284
		when 000645 => D <= "00000100";	-- 0x0285
		when 000646 => D <= "00100001";	-- 0x0286
		when 000647 => D <= "00000000";	-- 0x0287
		when 000648 => D <= "00000000";	-- 0x0288
		when 000649 => D <= "11001101";	-- 0x0289
		when 000650 => D <= "01111010";	-- 0x028A
		when 000651 => D <= "00100001";	-- 0x028B
		when 000652 => D <= "00001110";	-- 0x028C
		when 000653 => D <= "00001000";	-- 0x028D
		when 000654 => D <= "00111110";	-- 0x028E
		when 000655 => D <= "00001011";	-- 0x028F
		when 000656 => D <= "11001101";	-- 0x0290
		when 000657 => D <= "11110011";	-- 0x0291
		when 000658 => D <= "00100000";	-- 0x0292
		when 000659 => D <= "00001101";	-- 0x0293
		when 000660 => D <= "11000010";	-- 0x0294
		when 000661 => D <= "10001110";	-- 0x0295
		when 000662 => D <= "00100010";	-- 0x0296
		when 000663 => D <= "00100001";	-- 0x0297
		when 000664 => D <= "01000000";	-- 0x0298
		when 000665 => D <= "00000000";	-- 0x0299
		when 000666 => D <= "00011001";	-- 0x029A
		when 000667 => D <= "11101011";	-- 0x029B
		when 000668 => D <= "00000101";	-- 0x029C
		when 000669 => D <= "11000010";	-- 0x029D
		when 000670 => D <= "10000110";	-- 0x029E
		when 000671 => D <= "00100010";	-- 0x029F
		when 000672 => D <= "00111110";	-- 0x02A0
		when 000673 => D <= "00010001";	-- 0x02A1
		when 000674 => D <= "11000011";	-- 0x02A2
		when 000675 => D <= "01101000";	-- 0x02A3
		when 000676 => D <= "00100010";	-- 0x02A4
		when 000677 => D <= "00010001";	-- 0x02A5
		when 000678 => D <= "01101000";	-- 0x02A6
		when 000679 => D <= "00000001";	-- 0x02A7
		when 000680 => D <= "01111100";	-- 0x02A8
		when 000681 => D <= "10110111";	-- 0x02A9
		when 000682 => D <= "11111010";	-- 0x02AA
		when 000683 => D <= "11000001";	-- 0x02AB
		when 000684 => D <= "00100010";	-- 0x02AC
		when 000685 => D <= "11100101";	-- 0x02AD
		when 000686 => D <= "00100001";	-- 0x02AE
		when 000687 => D <= "10111110";	-- 0x02AF
		when 000688 => D <= "00100010";	-- 0x02B0
		when 000689 => D <= "11100011";	-- 0x02B1
		when 000690 => D <= "11100101";	-- 0x02B2
		when 000691 => D <= "10101111";	-- 0x02B3
		when 000692 => D <= "11101101";	-- 0x02B4
		when 000693 => D <= "01010010";	-- 0x02B5
		when 000694 => D <= "11100001";	-- 0x02B6
		when 000695 => D <= "11111000";	-- 0x02B7
		when 000696 => D <= "10101111";	-- 0x02B8
		when 000697 => D <= "11101101";	-- 0x02B9
		when 000698 => D <= "01010010";	-- 0x02BA
		when 000699 => D <= "11000011";	-- 0x02BB
		when 000700 => D <= "10110010";	-- 0x02BC
		when 000701 => D <= "00100010";	-- 0x02BD
		when 000702 => D <= "11000011";	-- 0x02BE
		when 000703 => D <= "11000111";	-- 0x02BF
		when 000704 => D <= "00100010";	-- 0x02C0
		when 000705 => D <= "00011001";	-- 0x02C1
		when 000706 => D <= "01111100";	-- 0x02C2
		when 000707 => D <= "10110111";	-- 0x02C3
		when 000708 => D <= "11111010";	-- 0x02C4
		when 000709 => D <= "11000001";	-- 0x02C5
		when 000710 => D <= "00100010";	-- 0x02C6
		when 000711 => D <= "11001001";	-- 0x02C7
		when 000712 => D <= "00001110";	-- 0x02C8
		when 000713 => D <= "00000000";	-- 0x02C9
		when 000714 => D <= "01111010";	-- 0x02CA
		when 000715 => D <= "10110111";	-- 0x02CB
		when 000716 => D <= "11110010";	-- 0x02CC
		when 000717 => D <= "11010111";	-- 0x02CD
		when 000718 => D <= "00100010";	-- 0x02CE
		when 000719 => D <= "00001110";	-- 0x02CF
		when 000720 => D <= "00000001";	-- 0x02D0
		when 000721 => D <= "00101111";	-- 0x02D1
		when 000722 => D <= "01010111";	-- 0x02D2
		when 000723 => D <= "01111011";	-- 0x02D3
		when 000724 => D <= "00101111";	-- 0x02D4
		when 000725 => D <= "01011111";	-- 0x02D5
		when 000726 => D <= "00010011";	-- 0x02D6
		when 000727 => D <= "01111000";	-- 0x02D7
		when 000728 => D <= "10101001";	-- 0x02D8
		when 000729 => D <= "00110010";	-- 0x02D9
		when 000730 => D <= "00101111";	-- 0x02DA
		when 000731 => D <= "10000000";	-- 0x02DB
		when 000732 => D <= "11001011";	-- 0x02DC
		when 000733 => D <= "01000100";	-- 0x02DD
		when 000734 => D <= "11000010";	-- 0x02DE
		when 000735 => D <= "00000010";	-- 0x02DF
		when 000736 => D <= "00100011";	-- 0x02E0
		when 000737 => D <= "01111101";	-- 0x02E1
		when 000738 => D <= "00001110";	-- 0x02E2
		when 000739 => D <= "00001000";	-- 0x02E3
		when 000740 => D <= "00100001";	-- 0x02E4
		when 000741 => D <= "00000000";	-- 0x02E5
		when 000742 => D <= "00000000";	-- 0x02E6
		when 000743 => D <= "00101001";	-- 0x02E7
		when 000744 => D <= "00010111";	-- 0x02E8
		when 000745 => D <= "11010010";	-- 0x02E9
		when 000746 => D <= "11101111";	-- 0x02EA
		when 000747 => D <= "00100010";	-- 0x02EB
		when 000748 => D <= "00011001";	-- 0x02EC
		when 000749 => D <= "11001110";	-- 0x02ED
		when 000750 => D <= "00000000";	-- 0x02EE
		when 000751 => D <= "00001101";	-- 0x02EF
		when 000752 => D <= "11000010";	-- 0x02F0
		when 000753 => D <= "11100111";	-- 0x02F1
		when 000754 => D <= "00100010";	-- 0x02F2
		when 000755 => D <= "01101100";	-- 0x02F3
		when 000756 => D <= "01100111";	-- 0x02F4
		when 000757 => D <= "00111010";	-- 0x02F5
		when 000758 => D <= "00101111";	-- 0x02F6
		when 000759 => D <= "10000000";	-- 0x02F7
		when 000760 => D <= "10110111";	-- 0x02F8
		when 000761 => D <= "11001000";	-- 0x02F9
		when 000762 => D <= "01111100";	-- 0x02FA
		when 000763 => D <= "00101111";	-- 0x02FB
		when 000764 => D <= "01100111";	-- 0x02FC
		when 000765 => D <= "01111101";	-- 0x02FD
		when 000766 => D <= "00101111";	-- 0x02FE
		when 000767 => D <= "01101111";	-- 0x02FF
		when 000768 => D <= "00100011";	-- 0x0300
		when 000769 => D <= "11001001";	-- 0x0301
		when 000770 => D <= "11101011";	-- 0x0302
		when 000771 => D <= "11000011";	-- 0x0303
		when 000772 => D <= "11110101";	-- 0x0304
		when 000773 => D <= "00100010";	-- 0x0305
		when 000774 => D <= "00000000";	-- 0x0306
		when 000775 => D <= "00000100";	-- 0x0307
		when 000776 => D <= "00001001";	-- 0x0308
		when 000777 => D <= "00001101";	-- 0x0309
		when 000778 => D <= "00010010";	-- 0x030A
		when 000779 => D <= "00010110";	-- 0x030B
		when 000780 => D <= "00011011";	-- 0x030C
		when 000781 => D <= "00011111";	-- 0x030D
		when 000782 => D <= "00100100";	-- 0x030E
		when 000783 => D <= "00101000";	-- 0x030F
		when 000784 => D <= "00101100";	-- 0x0310
		when 000785 => D <= "00110001";	-- 0x0311
		when 000786 => D <= "00110101";	-- 0x0312
		when 000787 => D <= "00111010";	-- 0x0313
		when 000788 => D <= "00111110";	-- 0x0314
		when 000789 => D <= "01000010";	-- 0x0315
		when 000790 => D <= "01000111";	-- 0x0316
		when 000791 => D <= "01001011";	-- 0x0317
		when 000792 => D <= "01001111";	-- 0x0318
		when 000793 => D <= "01010011";	-- 0x0319
		when 000794 => D <= "01011000";	-- 0x031A
		when 000795 => D <= "01011100";	-- 0x031B
		when 000796 => D <= "01100000";	-- 0x031C
		when 000797 => D <= "01100100";	-- 0x031D
		when 000798 => D <= "01101000";	-- 0x031E
		when 000799 => D <= "01101100";	-- 0x031F
		when 000800 => D <= "01110000";	-- 0x0320
		when 000801 => D <= "01110100";	-- 0x0321
		when 000802 => D <= "01111000";	-- 0x0322
		when 000803 => D <= "01111100";	-- 0x0323
		when 000804 => D <= "10000000";	-- 0x0324
		when 000805 => D <= "10000100";	-- 0x0325
		when 000806 => D <= "10001000";	-- 0x0326
		when 000807 => D <= "10001011";	-- 0x0327
		when 000808 => D <= "10001111";	-- 0x0328
		when 000809 => D <= "10010011";	-- 0x0329
		when 000810 => D <= "10010110";	-- 0x032A
		when 000811 => D <= "10011010";	-- 0x032B
		when 000812 => D <= "10011110";	-- 0x032C
		when 000813 => D <= "10100001";	-- 0x032D
		when 000814 => D <= "10100101";	-- 0x032E
		when 000815 => D <= "10101000";	-- 0x032F
		when 000816 => D <= "10101011";	-- 0x0330
		when 000817 => D <= "10101111";	-- 0x0331
		when 000818 => D <= "10110010";	-- 0x0332
		when 000819 => D <= "10110101";	-- 0x0333
		when 000820 => D <= "10111000";	-- 0x0334
		when 000821 => D <= "10111011";	-- 0x0335
		when 000822 => D <= "10111110";	-- 0x0336
		when 000823 => D <= "11000001";	-- 0x0337
		when 000824 => D <= "11000100";	-- 0x0338
		when 000825 => D <= "11000111";	-- 0x0339
		when 000826 => D <= "11001010";	-- 0x033A
		when 000827 => D <= "11001100";	-- 0x033B
		when 000828 => D <= "11001111";	-- 0x033C
		when 000829 => D <= "11010010";	-- 0x033D
		when 000830 => D <= "11010100";	-- 0x033E
		when 000831 => D <= "11010111";	-- 0x033F
		when 000832 => D <= "11011001";	-- 0x0340
		when 000833 => D <= "11011011";	-- 0x0341
		when 000834 => D <= "11011110";	-- 0x0342
		when 000835 => D <= "11100000";	-- 0x0343
		when 000836 => D <= "11100010";	-- 0x0344
		when 000837 => D <= "11100100";	-- 0x0345
		when 000838 => D <= "11100110";	-- 0x0346
		when 000839 => D <= "11101000";	-- 0x0347
		when 000840 => D <= "11101010";	-- 0x0348
		when 000841 => D <= "11101100";	-- 0x0349
		when 000842 => D <= "11101101";	-- 0x034A
		when 000843 => D <= "11101111";	-- 0x034B
		when 000844 => D <= "11110001";	-- 0x034C
		when 000845 => D <= "11110010";	-- 0x034D
		when 000846 => D <= "11110011";	-- 0x034E
		when 000847 => D <= "11110101";	-- 0x034F
		when 000848 => D <= "11110110";	-- 0x0350
		when 000849 => D <= "11110111";	-- 0x0351
		when 000850 => D <= "11111000";	-- 0x0352
		when 000851 => D <= "11111001";	-- 0x0353
		when 000852 => D <= "11111010";	-- 0x0354
		when 000853 => D <= "11111011";	-- 0x0355
		when 000854 => D <= "11111100";	-- 0x0356
		when 000855 => D <= "11111101";	-- 0x0357
		when 000856 => D <= "11111110";	-- 0x0358
		when 000857 => D <= "11111110";	-- 0x0359
		when 000858 => D <= "11111111";	-- 0x035A
		when 000859 => D <= "11111111";	-- 0x035B
		when 000860 => D <= "11111111";	-- 0x035C
		when 000861 => D <= "00000000";	-- 0x035D
		when 000862 => D <= "00000000";	-- 0x035E
		when 000863 => D <= "00000000";	-- 0x035F
		when 000864 => D <= "00000000";	-- 0x0360
		when 000865 => D <= "11101011";	-- 0x0361
		when 000866 => D <= "00100001";	-- 0x0362
		when 000867 => D <= "01011010";	-- 0x0363
		when 000868 => D <= "00000000";	-- 0x0364
		when 000869 => D <= "10101111";	-- 0x0365
		when 000870 => D <= "11101101";	-- 0x0366
		when 000871 => D <= "01010010";	-- 0x0367
		when 000872 => D <= "11001011";	-- 0x0368
		when 000873 => D <= "01111100";	-- 0x0369
		when 000874 => D <= "11001010";	-- 0x036A
		when 000875 => D <= "01110001";	-- 0x036B
		when 000876 => D <= "00100011";	-- 0x036C
		when 000877 => D <= "00010001";	-- 0x036D
		when 000878 => D <= "01101000";	-- 0x036E
		when 000879 => D <= "00000001";	-- 0x036F
		when 000880 => D <= "00011001";	-- 0x0370
		when 000881 => D <= "00100010";	-- 0x0371
		when 000882 => D <= "00110100";	-- 0x0372
		when 000883 => D <= "10000000";	-- 0x0373
		when 000884 => D <= "00000110";	-- 0x0374
		when 000885 => D <= "00000000";	-- 0x0375
		when 000886 => D <= "00010001";	-- 0x0376
		when 000887 => D <= "01011010";	-- 0x0377
		when 000888 => D <= "00000000";	-- 0x0378
		when 000889 => D <= "10101111";	-- 0x0379
		when 000890 => D <= "11101101";	-- 0x037A
		when 000891 => D <= "01010010";	-- 0x037B
		when 000892 => D <= "11111010";	-- 0x037C
		when 000893 => D <= "10111001";	-- 0x037D
		when 000894 => D <= "00100011";	-- 0x037E
		when 000895 => D <= "00010001";	-- 0x037F
		when 000896 => D <= "01011010";	-- 0x0380
		when 000897 => D <= "00000000";	-- 0x0381
		when 000898 => D <= "10101111";	-- 0x0382
		when 000899 => D <= "11101101";	-- 0x0383
		when 000900 => D <= "01010010";	-- 0x0384
		when 000901 => D <= "11111010";	-- 0x0385
		when 000902 => D <= "10101100";	-- 0x0386
		when 000903 => D <= "00100011";	-- 0x0387
		when 000904 => D <= "00000110";	-- 0x0388
		when 000905 => D <= "00000001";	-- 0x0389
		when 000906 => D <= "00010001";	-- 0x038A
		when 000907 => D <= "01011010";	-- 0x038B
		when 000908 => D <= "00000000";	-- 0x038C
		when 000909 => D <= "10101111";	-- 0x038D
		when 000910 => D <= "11101101";	-- 0x038E
		when 000911 => D <= "01010010";	-- 0x038F
		when 000912 => D <= "11111010";	-- 0x0390
		when 000913 => D <= "10100000";	-- 0x0391
		when 000914 => D <= "00100011";	-- 0x0392
		when 000915 => D <= "00100001";	-- 0x0393
		when 000916 => D <= "01101000";	-- 0x0394
		when 000917 => D <= "00000001";	-- 0x0395
		when 000918 => D <= "11101101";	-- 0x0396
		when 000919 => D <= "01011011";	-- 0x0397
		when 000920 => D <= "00110100";	-- 0x0398
		when 000921 => D <= "10000000";	-- 0x0399
		when 000922 => D <= "10101111";	-- 0x039A
		when 000923 => D <= "11101101";	-- 0x039B
		when 000924 => D <= "01010010";	-- 0x039C
		when 000925 => D <= "11000011";	-- 0x039D
		when 000926 => D <= "10101001";	-- 0x039E
		when 000927 => D <= "00100011";	-- 0x039F
		when 000928 => D <= "00101010";	-- 0x03A0
		when 000929 => D <= "00110100";	-- 0x03A1
		when 000930 => D <= "10000000";	-- 0x03A2
		when 000931 => D <= "00010001";	-- 0x03A3
		when 000932 => D <= "10110100";	-- 0x03A4
		when 000933 => D <= "00000000";	-- 0x03A5
		when 000934 => D <= "10101111";	-- 0x03A6
		when 000935 => D <= "11101101";	-- 0x03A7
		when 000936 => D <= "01010010";	-- 0x03A8
		when 000937 => D <= "11000011";	-- 0x03A9
		when 000938 => D <= "10110110";	-- 0x03AA
		when 000939 => D <= "00100011";	-- 0x03AB
		when 000940 => D <= "11101101";	-- 0x03AC
		when 000941 => D <= "01011011";	-- 0x03AD
		when 000942 => D <= "00110100";	-- 0x03AE
		when 000943 => D <= "10000000";	-- 0x03AF
		when 000944 => D <= "00100001";	-- 0x03B0
		when 000945 => D <= "10110100";	-- 0x03B1
		when 000946 => D <= "00000000";	-- 0x03B2
		when 000947 => D <= "10101111";	-- 0x03B3
		when 000948 => D <= "11101101";	-- 0x03B4
		when 000949 => D <= "01010010";	-- 0x03B5
		when 000950 => D <= "11000011";	-- 0x03B6
		when 000951 => D <= "10111100";	-- 0x03B7
		when 000952 => D <= "00100011";	-- 0x03B8
		when 000953 => D <= "00101010";	-- 0x03B9
		when 000954 => D <= "00110100";	-- 0x03BA
		when 000955 => D <= "10000000";	-- 0x03BB
		when 000956 => D <= "01111100";	-- 0x03BC
		when 000957 => D <= "10110101";	-- 0x03BD
		when 000958 => D <= "11001000";	-- 0x03BE
		when 000959 => D <= "11101011";	-- 0x03BF
		when 000960 => D <= "00100001";	-- 0x03C0
		when 000961 => D <= "00000110";	-- 0x03C1
		when 000962 => D <= "00100011";	-- 0x03C2
		when 000963 => D <= "00011001";	-- 0x03C3
		when 000964 => D <= "01101110";	-- 0x03C4
		when 000965 => D <= "00100110";	-- 0x03C5
		when 000966 => D <= "00000000";	-- 0x03C6
		when 000967 => D <= "01111101";	-- 0x03C7
		when 000968 => D <= "10110111";	-- 0x03C8
		when 000969 => D <= "11000000";	-- 0x03C9
		when 000970 => D <= "00100110";	-- 0x03CA
		when 000971 => D <= "00000001";	-- 0x03CB
		when 000972 => D <= "11001001";	-- 0x03CC
		when 000973 => D <= "11001101";	-- 0x03CD
		when 000974 => D <= "11101010";	-- 0x03CE
		when 000975 => D <= "00100000";	-- 0x03CF
		when 000976 => D <= "11011011";	-- 0x03D0
		when 000977 => D <= "01111000";	-- 0x03D1
		when 000978 => D <= "00110010";	-- 0x03D2
		when 000979 => D <= "00110001";	-- 0x03D3
		when 000980 => D <= "10000000";	-- 0x03D4
		when 000981 => D <= "11011011";	-- 0x03D5
		when 000982 => D <= "01111001";	-- 0x03D6
		when 000983 => D <= "00110010";	-- 0x03D7
		when 000984 => D <= "00110000";	-- 0x03D8
		when 000985 => D <= "10000000";	-- 0x03D9
		when 000986 => D <= "11011011";	-- 0x03DA
		when 000987 => D <= "01111010";	-- 0x03DB
		when 000988 => D <= "00110010";	-- 0x03DC
		when 000989 => D <= "00110011";	-- 0x03DD
		when 000990 => D <= "10000000";	-- 0x03DE
		when 000991 => D <= "11011011";	-- 0x03DF
		when 000992 => D <= "01111011";	-- 0x03E0
		when 000993 => D <= "00110010";	-- 0x03E1
		when 000994 => D <= "00110010";	-- 0x03E2
		when 000995 => D <= "10000000";	-- 0x03E3
		when 000996 => D <= "11001001";	-- 0x03E4
		when 000997 => D <= "11001101";	-- 0x03E5
		when 000998 => D <= "11101010";	-- 0x03E6
		when 000999 => D <= "00100000";	-- 0x03E7
		when 001000 => D <= "00111010";	-- 0x03E8
		when 001001 => D <= "00110001";	-- 0x03E9
		when 001002 => D <= "10000000";	-- 0x03EA
		when 001003 => D <= "11010011";	-- 0x03EB
		when 001004 => D <= "01111000";	-- 0x03EC
		when 001005 => D <= "00111010";	-- 0x03ED
		when 001006 => D <= "00110000";	-- 0x03EE
		when 001007 => D <= "10000000";	-- 0x03EF
		when 001008 => D <= "11010011";	-- 0x03F0
		when 001009 => D <= "01111001";	-- 0x03F1
		when 001010 => D <= "00111010";	-- 0x03F2
		when 001011 => D <= "00110011";	-- 0x03F3
		when 001012 => D <= "10000000";	-- 0x03F4
		when 001013 => D <= "11010011";	-- 0x03F5
		when 001014 => D <= "01111010";	-- 0x03F6
		when 001015 => D <= "00111010";	-- 0x03F7
		when 001016 => D <= "00110010";	-- 0x03F8
		when 001017 => D <= "10000000";	-- 0x03F9
		when 001018 => D <= "11010011";	-- 0x03FA
		when 001019 => D <= "01111011";	-- 0x03FB
		when 001020 => D <= "11001001";	-- 0x03FC
		when 001021 => D <= "00100001";	-- 0x03FD
		when 001022 => D <= "00000000";	-- 0x03FE
		when 001023 => D <= "00000001";	-- 0x03FF
		when 001024 => D <= "00010001";	-- 0x0400
		when 001025 => D <= "00000000";	-- 0x0401
		when 001026 => D <= "00000001";	-- 0x0402
		when 001027 => D <= "00000001";	-- 0x0403
		when 001028 => D <= "01011010";	-- 0x0404
		when 001029 => D <= "00000000";	-- 0x0405
		when 001030 => D <= "11000011";	-- 0x0406
		when 001031 => D <= "00001001";	-- 0x0407
		when 001032 => D <= "00100100";	-- 0x0408
		when 001033 => D <= "11001101";	-- 0x0409
		when 001034 => D <= "00010100";	-- 0x040A
		when 001035 => D <= "00100101";	-- 0x040B
		when 001036 => D <= "00100010";	-- 0x040C
		when 001037 => D <= "00110111";	-- 0x040D
		when 001038 => D <= "10000000";	-- 0x040E
		when 001039 => D <= "11101011";	-- 0x040F
		when 001040 => D <= "11001101";	-- 0x0410
		when 001041 => D <= "00010100";	-- 0x0411
		when 001042 => D <= "00100101";	-- 0x0412
		when 001043 => D <= "00100010";	-- 0x0413
		when 001044 => D <= "00111001";	-- 0x0414
		when 001045 => D <= "10000000";	-- 0x0415
		when 001046 => D <= "01101001";	-- 0x0416
		when 001047 => D <= "01100000";	-- 0x0417
		when 001048 => D <= "11001101";	-- 0x0418
		when 001049 => D <= "10100101";	-- 0x0419
		when 001050 => D <= "00100010";	-- 0x041A
		when 001051 => D <= "00100010";	-- 0x041B
		when 001052 => D <= "00111011";	-- 0x041C
		when 001053 => D <= "10000000";	-- 0x041D
		when 001054 => D <= "11001101";	-- 0x041E
		when 001055 => D <= "00011110";	-- 0x041F
		when 001056 => D <= "00100101";	-- 0x0420
		when 001057 => D <= "00111110";	-- 0x0421
		when 001058 => D <= "00000001";	-- 0x0422
		when 001059 => D <= "00110010";	-- 0x0423
		when 001060 => D <= "00100111";	-- 0x0424
		when 001061 => D <= "10000000";	-- 0x0425
		when 001062 => D <= "00110010";	-- 0x0426
		when 001063 => D <= "00101000";	-- 0x0427
		when 001064 => D <= "10000000";	-- 0x0428
		when 001065 => D <= "10101111";	-- 0x0429
		when 001066 => D <= "00110010";	-- 0x042A
		when 001067 => D <= "00110110";	-- 0x042B
		when 001068 => D <= "10000000";	-- 0x042C
		when 001069 => D <= "11001001";	-- 0x042D
		when 001070 => D <= "00111010";	-- 0x042E
		when 001071 => D <= "00110110";	-- 0x042F
		when 001072 => D <= "10000000";	-- 0x0430
		when 001073 => D <= "11111110";	-- 0x0431
		when 001074 => D <= "00000001";	-- 0x0432
		when 001075 => D <= "11000010";	-- 0x0433
		when 001076 => D <= "00111001";	-- 0x0434
		when 001077 => D <= "00100100";	-- 0x0435
		when 001078 => D <= "11001101";	-- 0x0436
		when 001079 => D <= "11111101";	-- 0x0437
		when 001080 => D <= "00100011";	-- 0x0438
		when 001081 => D <= "11001001";	-- 0x0439
		when 001082 => D <= "11011101";	-- 0x043A
		when 001083 => D <= "11100101";	-- 0x043B
		when 001084 => D <= "11001101";	-- 0x043C
		when 001085 => D <= "00101110";	-- 0x043D
		when 001086 => D <= "00100100";	-- 0x043E
		when 001087 => D <= "00111010";	-- 0x043F
		when 001088 => D <= "01000111";	-- 0x0440
		when 001089 => D <= "10000000";	-- 0x0441
		when 001090 => D <= "00110010";	-- 0x0442
		when 001091 => D <= "01000110";	-- 0x0443
		when 001092 => D <= "10000000";	-- 0x0444
		when 001093 => D <= "11001101";	-- 0x0445
		when 001094 => D <= "01011000";	-- 0x0446
		when 001095 => D <= "00100001";	-- 0x0447
		when 001096 => D <= "00111010";	-- 0x0448
		when 001097 => D <= "00101001";	-- 0x0449
		when 001098 => D <= "10000000";	-- 0x044A
		when 001099 => D <= "11001101";	-- 0x044B
		when 001100 => D <= "11110011";	-- 0x044C
		when 001101 => D <= "00100000";	-- 0x044D
		when 001102 => D <= "00101010";	-- 0x044E
		when 001103 => D <= "00110111";	-- 0x044F
		when 001104 => D <= "10000000";	-- 0x0450
		when 001105 => D <= "11101101";	-- 0x0451
		when 001106 => D <= "01011011";	-- 0x0452
		when 001107 => D <= "00111001";	-- 0x0453
		when 001108 => D <= "10000000";	-- 0x0454
		when 001109 => D <= "11001101";	-- 0x0455
		when 001110 => D <= "11011010";	-- 0x0456
		when 001111 => D <= "00100101";	-- 0x0457
		when 001112 => D <= "11001101";	-- 0x0458
		when 001113 => D <= "01111010";	-- 0x0459
		when 001114 => D <= "00100001";	-- 0x045A
		when 001115 => D <= "11011101";	-- 0x045B
		when 001116 => D <= "11100001";	-- 0x045C
		when 001117 => D <= "11001001";	-- 0x045D
		when 001118 => D <= "11001101";	-- 0x045E
		when 001119 => D <= "00010100";	-- 0x045F
		when 001120 => D <= "00100101";	-- 0x0460
		when 001121 => D <= "11110101";	-- 0x0461
		when 001122 => D <= "11000101";	-- 0x0462
		when 001123 => D <= "11010101";	-- 0x0463
		when 001124 => D <= "11100101";	-- 0x0464
		when 001125 => D <= "11100101";	-- 0x0465
		when 001126 => D <= "11001101";	-- 0x0466
		when 001127 => D <= "00111010";	-- 0x0467
		when 001128 => D <= "00100100";	-- 0x0468
		when 001129 => D <= "00101010";	-- 0x0469
		when 001130 => D <= "00111011";	-- 0x046A
		when 001131 => D <= "10000000";	-- 0x046B
		when 001132 => D <= "11001101";	-- 0x046C
		when 001133 => D <= "01100001";	-- 0x046D
		when 001134 => D <= "00100011";	-- 0x046E
		when 001135 => D <= "11010001";	-- 0x046F
		when 001136 => D <= "11010101";	-- 0x0470
		when 001137 => D <= "11001101";	-- 0x0471
		when 001138 => D <= "11001000";	-- 0x0472
		when 001139 => D <= "00100010";	-- 0x0473
		when 001140 => D <= "11101101";	-- 0x0474
		when 001141 => D <= "01011011";	-- 0x0475
		when 001142 => D <= "00110111";	-- 0x0476
		when 001143 => D <= "10000000";	-- 0x0477
		when 001144 => D <= "00011001";	-- 0x0478
		when 001145 => D <= "00100010";	-- 0x0479
		when 001146 => D <= "00110111";	-- 0x047A
		when 001147 => D <= "10000000";	-- 0x047B
		when 001148 => D <= "00101010";	-- 0x047C
		when 001149 => D <= "00111011";	-- 0x047D
		when 001150 => D <= "10000000";	-- 0x047E
		when 001151 => D <= "11001101";	-- 0x047F
		when 001152 => D <= "01110001";	-- 0x0480
		when 001153 => D <= "00100011";	-- 0x0481
		when 001154 => D <= "11010001";	-- 0x0482
		when 001155 => D <= "11001101";	-- 0x0483
		when 001156 => D <= "11001000";	-- 0x0484
		when 001157 => D <= "00100010";	-- 0x0485
		when 001158 => D <= "11101101";	-- 0x0486
		when 001159 => D <= "01011011";	-- 0x0487
		when 001160 => D <= "00111001";	-- 0x0488
		when 001161 => D <= "10000000";	-- 0x0489
		when 001162 => D <= "00011001";	-- 0x048A
		when 001163 => D <= "00100010";	-- 0x048B
		when 001164 => D <= "00111001";	-- 0x048C
		when 001165 => D <= "10000000";	-- 0x048D
		when 001166 => D <= "11001101";	-- 0x048E
		when 001167 => D <= "10010011";	-- 0x048F
		when 001168 => D <= "00100100";	-- 0x0490
		when 001169 => D <= "00011000";	-- 0x0491
		when 001170 => D <= "00110000";	-- 0x0492
		when 001171 => D <= "00101010";	-- 0x0493
		when 001172 => D <= "00110111";	-- 0x0494
		when 001173 => D <= "10000000";	-- 0x0495
		when 001174 => D <= "11101101";	-- 0x0496
		when 001175 => D <= "01011011";	-- 0x0497
		when 001176 => D <= "00111001";	-- 0x0498
		when 001177 => D <= "10000000";	-- 0x0499
		when 001178 => D <= "11001101";	-- 0x049A
		when 001179 => D <= "11011010";	-- 0x049B
		when 001180 => D <= "00100101";	-- 0x049C
		when 001181 => D <= "00111010";	-- 0x049D
		when 001182 => D <= "01000011";	-- 0x049E
		when 001183 => D <= "10000000";	-- 0x049F
		when 001184 => D <= "11111110";	-- 0x04A0
		when 001185 => D <= "00000001";	-- 0x04A1
		when 001186 => D <= "11000010";	-- 0x04A2
		when 001187 => D <= "10101011";	-- 0x04A3
		when 001188 => D <= "00100100";	-- 0x04A4
		when 001189 => D <= "11001101";	-- 0x04A5
		when 001190 => D <= "10001010";	-- 0x04A6
		when 001191 => D <= "00100001";	-- 0x04A7
		when 001192 => D <= "11000011";	-- 0x04A8
		when 001193 => D <= "10101110";	-- 0x04A9
		when 001194 => D <= "00100100";	-- 0x04AA
		when 001195 => D <= "11001101";	-- 0x04AB
		when 001196 => D <= "01111010";	-- 0x04AC
		when 001197 => D <= "00100001";	-- 0x04AD
		when 001198 => D <= "11001001";	-- 0x04AE
		when 001199 => D <= "11110101";	-- 0x04AF
		when 001200 => D <= "11000101";	-- 0x04B0
		when 001201 => D <= "11010101";	-- 0x04B1
		when 001202 => D <= "11100101";	-- 0x04B2
		when 001203 => D <= "11100101";	-- 0x04B3
		when 001204 => D <= "11001101";	-- 0x04B4
		when 001205 => D <= "00101110";	-- 0x04B5
		when 001206 => D <= "00100100";	-- 0x04B6
		when 001207 => D <= "11100001";	-- 0x04B7
		when 001208 => D <= "11101101";	-- 0x04B8
		when 001209 => D <= "01011011";	-- 0x04B9
		when 001210 => D <= "00111011";	-- 0x04BA
		when 001211 => D <= "10000000";	-- 0x04BB
		when 001212 => D <= "00011001";	-- 0x04BC
		when 001213 => D <= "11001101";	-- 0x04BD
		when 001214 => D <= "10100101";	-- 0x04BE
		when 001215 => D <= "00100010";	-- 0x04BF
		when 001216 => D <= "00100010";	-- 0x04C0
		when 001217 => D <= "00111011";	-- 0x04C1
		when 001218 => D <= "10000000";	-- 0x04C2
		when 001219 => D <= "11001101";	-- 0x04C3
		when 001220 => D <= "01011001";	-- 0x04C4
		when 001221 => D <= "00100000";	-- 0x04C5
		when 001222 => D <= "11100001";	-- 0x04C6
		when 001223 => D <= "11010001";	-- 0x04C7
		when 001224 => D <= "11000001";	-- 0x04C8
		when 001225 => D <= "11110001";	-- 0x04C9
		when 001226 => D <= "11001001";	-- 0x04CA
		when 001227 => D <= "11110101";	-- 0x04CB
		when 001228 => D <= "10101111";	-- 0x04CC
		when 001229 => D <= "00110010";	-- 0x04CD
		when 001230 => D <= "01000011";	-- 0x04CE
		when 001231 => D <= "10000000";	-- 0x04CF
		when 001232 => D <= "11110001";	-- 0x04D0
		when 001233 => D <= "11001001";	-- 0x04D1
		when 001234 => D <= "11110101";	-- 0x04D2
		when 001235 => D <= "00111110";	-- 0x04D3
		when 001236 => D <= "00000001";	-- 0x04D4
		when 001237 => D <= "00110010";	-- 0x04D5
		when 001238 => D <= "01000011";	-- 0x04D6
		when 001239 => D <= "10000000";	-- 0x04D7
		when 001240 => D <= "11110001";	-- 0x04D8
		when 001241 => D <= "11001001";	-- 0x04D9
		when 001242 => D <= "00111010";	-- 0x04DA
		when 001243 => D <= "00110110";	-- 0x04DB
		when 001244 => D <= "10000000";	-- 0x04DC
		when 001245 => D <= "11111110";	-- 0x04DD
		when 001246 => D <= "00000001";	-- 0x04DE
		when 001247 => D <= "11000010";	-- 0x04DF
		when 001248 => D <= "11100101";	-- 0x04E0
		when 001249 => D <= "00100100";	-- 0x04E1
		when 001250 => D <= "11001101";	-- 0x04E2
		when 001251 => D <= "11111101";	-- 0x04E3
		when 001252 => D <= "00100011";	-- 0x04E4
		when 001253 => D <= "10101111";	-- 0x04E5
		when 001254 => D <= "00110010";	-- 0x04E6
		when 001255 => D <= "00100111";	-- 0x04E7
		when 001256 => D <= "10000000";	-- 0x04E8
		when 001257 => D <= "00110010";	-- 0x04E9
		when 001258 => D <= "00100101";	-- 0x04EA
		when 001259 => D <= "10000000";	-- 0x04EB
		when 001260 => D <= "00110010";	-- 0x04EC
		when 001261 => D <= "01000101";	-- 0x04ED
		when 001262 => D <= "10000000";	-- 0x04EE
		when 001263 => D <= "00110010";	-- 0x04EF
		when 001264 => D <= "01000110";	-- 0x04F0
		when 001265 => D <= "10000000";	-- 0x04F1
		when 001266 => D <= "11001101";	-- 0x04F2
		when 001267 => D <= "01011000";	-- 0x04F3
		when 001268 => D <= "00100001";	-- 0x04F4
		when 001269 => D <= "11001001";	-- 0x04F5
		when 001270 => D <= "00111010";	-- 0x04F6
		when 001271 => D <= "00110110";	-- 0x04F7
		when 001272 => D <= "10000000";	-- 0x04F8
		when 001273 => D <= "11111110";	-- 0x04F9
		when 001274 => D <= "00000001";	-- 0x04FA
		when 001275 => D <= "11000010";	-- 0x04FB
		when 001276 => D <= "00000001";	-- 0x04FC
		when 001277 => D <= "00100101";	-- 0x04FD
		when 001278 => D <= "11001101";	-- 0x04FE
		when 001279 => D <= "11111101";	-- 0x04FF
		when 001280 => D <= "00100011";	-- 0x0500
		when 001281 => D <= "00111110";	-- 0x0501
		when 001282 => D <= "00000001";	-- 0x0502
		when 001283 => D <= "00110010";	-- 0x0503
		when 001284 => D <= "00100111";	-- 0x0504
		when 001285 => D <= "10000000";	-- 0x0505
		when 001286 => D <= "00110010";	-- 0x0506
		when 001287 => D <= "00101000";	-- 0x0507
		when 001288 => D <= "10000000";	-- 0x0508
		when 001289 => D <= "10101111";	-- 0x0509
		when 001290 => D <= "00110010";	-- 0x050A
		when 001291 => D <= "01000101";	-- 0x050B
		when 001292 => D <= "10000000";	-- 0x050C
		when 001293 => D <= "00110010";	-- 0x050D
		when 001294 => D <= "01000110";	-- 0x050E
		when 001295 => D <= "10000000";	-- 0x050F
		when 001296 => D <= "11001101";	-- 0x0510
		when 001297 => D <= "01011000";	-- 0x0511
		when 001298 => D <= "00100001";	-- 0x0512
		when 001299 => D <= "11001001";	-- 0x0513
		when 001300 => D <= "00101001";	-- 0x0514
		when 001301 => D <= "00101001";	-- 0x0515
		when 001302 => D <= "00101001";	-- 0x0516
		when 001303 => D <= "00101001";	-- 0x0517
		when 001304 => D <= "11001001";	-- 0x0518
		when 001305 => D <= "00111010";	-- 0x0519
		when 001306 => D <= "00110110";	-- 0x051A
		when 001307 => D <= "10000000";	-- 0x051B
		when 001308 => D <= "10110111";	-- 0x051C
		when 001309 => D <= "11000000";	-- 0x051D
		when 001310 => D <= "11100101";	-- 0x051E
		when 001311 => D <= "11010101";	-- 0x051F
		when 001312 => D <= "11000101";	-- 0x0520
		when 001313 => D <= "00101010";	-- 0x0521
		when 001314 => D <= "00111101";	-- 0x0522
		when 001315 => D <= "10000000";	-- 0x0523
		when 001316 => D <= "11101101";	-- 0x0524
		when 001317 => D <= "01011011";	-- 0x0525
		when 001318 => D <= "00111111";	-- 0x0526
		when 001319 => D <= "10000000";	-- 0x0527
		when 001320 => D <= "11001101";	-- 0x0528
		when 001321 => D <= "11011010";	-- 0x0529
		when 001322 => D <= "00100101";	-- 0x052A
		when 001323 => D <= "11001101";	-- 0x052B
		when 001324 => D <= "01111010";	-- 0x052C
		when 001325 => D <= "00100001";	-- 0x052D
		when 001326 => D <= "00111110";	-- 0x052E
		when 001327 => D <= "00000001";	-- 0x052F
		when 001328 => D <= "00110010";	-- 0x0530
		when 001329 => D <= "01000110";	-- 0x0531
		when 001330 => D <= "10000000";	-- 0x0532
		when 001331 => D <= "11001101";	-- 0x0533
		when 001332 => D <= "01011000";	-- 0x0534
		when 001333 => D <= "00100001";	-- 0x0535
		when 001334 => D <= "11001101";	-- 0x0536
		when 001335 => D <= "01000110";	-- 0x0537
		when 001336 => D <= "00100010";	-- 0x0538
		when 001337 => D <= "11001101";	-- 0x0539
		when 001338 => D <= "01100111";	-- 0x053A
		when 001339 => D <= "00100101";	-- 0x053B
		when 001340 => D <= "00101010";	-- 0x053C
		when 001341 => D <= "00111011";	-- 0x053D
		when 001342 => D <= "10000000";	-- 0x053E
		when 001343 => D <= "00100010";	-- 0x053F
		when 001344 => D <= "01000001";	-- 0x0540
		when 001345 => D <= "10000000";	-- 0x0541
		when 001346 => D <= "00101010";	-- 0x0542
		when 001347 => D <= "00110111";	-- 0x0543
		when 001348 => D <= "10000000";	-- 0x0544
		when 001349 => D <= "00100010";	-- 0x0545
		when 001350 => D <= "00111101";	-- 0x0546
		when 001351 => D <= "10000000";	-- 0x0547
		when 001352 => D <= "11101101";	-- 0x0548
		when 001353 => D <= "01011011";	-- 0x0549
		when 001354 => D <= "00111001";	-- 0x054A
		when 001355 => D <= "10000000";	-- 0x054B
		when 001356 => D <= "11101101";	-- 0x054C
		when 001357 => D <= "01010011";	-- 0x054D
		when 001358 => D <= "00111111";	-- 0x054E
		when 001359 => D <= "10000000";	-- 0x054F
		when 001360 => D <= "11001101";	-- 0x0550
		when 001361 => D <= "11011010";	-- 0x0551
		when 001362 => D <= "00100101";	-- 0x0552
		when 001363 => D <= "11001101";	-- 0x0553
		when 001364 => D <= "01111010";	-- 0x0554
		when 001365 => D <= "00100001";	-- 0x0555
		when 001366 => D <= "11001101";	-- 0x0556
		when 001367 => D <= "01000010";	-- 0x0557
		when 001368 => D <= "00100010";	-- 0x0558
		when 001369 => D <= "11001101";	-- 0x0559
		when 001370 => D <= "01100111";	-- 0x055A
		when 001371 => D <= "00100101";	-- 0x055B
		when 001372 => D <= "10101111";	-- 0x055C
		when 001373 => D <= "00110010";	-- 0x055D
		when 001374 => D <= "01000110";	-- 0x055E
		when 001375 => D <= "10000000";	-- 0x055F
		when 001376 => D <= "11001101";	-- 0x0560
		when 001377 => D <= "01011000";	-- 0x0561
		when 001378 => D <= "00100001";	-- 0x0562
		when 001379 => D <= "11000001";	-- 0x0563
		when 001380 => D <= "11010001";	-- 0x0564
		when 001381 => D <= "11100001";	-- 0x0565
		when 001382 => D <= "11001001";	-- 0x0566
		when 001383 => D <= "00101010";	-- 0x0567
		when 001384 => D <= "01000001";	-- 0x0568
		when 001385 => D <= "10000000";	-- 0x0569
		when 001386 => D <= "10101111";	-- 0x056A
		when 001387 => D <= "00000110";	-- 0x056B
		when 001388 => D <= "00010000";	-- 0x056C
		when 001389 => D <= "11001011";	-- 0x056D
		when 001390 => D <= "00100101";	-- 0x056E
		when 001391 => D <= "11001011";	-- 0x056F
		when 001392 => D <= "00010100";	-- 0x0570
		when 001393 => D <= "00010111";	-- 0x0571
		when 001394 => D <= "11111110";	-- 0x0572
		when 001395 => D <= "00101101";	-- 0x0573
		when 001396 => D <= "11011010";	-- 0x0574
		when 001397 => D <= "01111011";	-- 0x0575
		when 001398 => D <= "00100101";	-- 0x0576
		when 001399 => D <= "11001011";	-- 0x0577
		when 001400 => D <= "11000101";	-- 0x0578
		when 001401 => D <= "11010110";	-- 0x0579
		when 001402 => D <= "00101101";	-- 0x057A
		when 001403 => D <= "00010000";	-- 0x057B
		when 001404 => D <= "11110000";	-- 0x057C
		when 001405 => D <= "00100110";	-- 0x057D
		when 001406 => D <= "00000000";	-- 0x057E
		when 001407 => D <= "01111101";	-- 0x057F
		when 001408 => D <= "11100110";	-- 0x0580
		when 001409 => D <= "00000111";	-- 0x0581
		when 001410 => D <= "01101111";	-- 0x0582
		when 001411 => D <= "00101001";	-- 0x0583
		when 001412 => D <= "00101001";	-- 0x0584
		when 001413 => D <= "00101001";	-- 0x0585
		when 001414 => D <= "00010001";	-- 0x0586
		when 001415 => D <= "10011010";	-- 0x0587
		when 001416 => D <= "00100101";	-- 0x0588
		when 001417 => D <= "00011001";	-- 0x0589
		when 001418 => D <= "00011110";	-- 0x058A
		when 001419 => D <= "00001000";	-- 0x058B
		when 001420 => D <= "01111110";	-- 0x058C
		when 001421 => D <= "10110111";	-- 0x058D
		when 001422 => D <= "11001010";	-- 0x058E
		when 001423 => D <= "10010100";	-- 0x058F
		when 001424 => D <= "00100101";	-- 0x0590
		when 001425 => D <= "11001101";	-- 0x0591
		when 001426 => D <= "11110011";	-- 0x0592
		when 001427 => D <= "00100000";	-- 0x0593
		when 001428 => D <= "00100011";	-- 0x0594
		when 001429 => D <= "00011101";	-- 0x0595
		when 001430 => D <= "11000010";	-- 0x0596
		when 001431 => D <= "10001100";	-- 0x0597
		when 001432 => D <= "00100101";	-- 0x0598
		when 001433 => D <= "11001001";	-- 0x0599
		when 001434 => D <= "11111010";	-- 0x059A
		when 001435 => D <= "11111101";	-- 0x059B
		when 001436 => D <= "11111111";	-- 0x059C
		when 001437 => D <= "11111010";	-- 0x059D
		when 001438 => D <= "00000000";	-- 0x059E
		when 001439 => D <= "00000000";	-- 0x059F
		when 001440 => D <= "00000000";	-- 0x05A0
		when 001441 => D <= "00000000";	-- 0x05A1
		when 001442 => D <= "11010011";	-- 0x05A2
		when 001443 => D <= "11010000";	-- 0x05A3
		when 001444 => D <= "11010000";	-- 0x05A4
		when 001445 => D <= "11010100";	-- 0x05A5
		when 001446 => D <= "11010100";	-- 0x05A6
		when 001447 => D <= "11010011";	-- 0x05A7
		when 001448 => D <= "00000000";	-- 0x05A8
		when 001449 => D <= "00000000";	-- 0x05A9
		when 001450 => D <= "11111110";	-- 0x05AA
		when 001451 => D <= "11111001";	-- 0x05AB
		when 001452 => D <= "11111101";	-- 0x05AC
		when 001453 => D <= "11111110";	-- 0x05AD
		when 001454 => D <= "00000000";	-- 0x05AE
		when 001455 => D <= "00000000";	-- 0x05AF
		when 001456 => D <= "00000000";	-- 0x05B0
		when 001457 => D <= "00000000";	-- 0x05B1
		when 001458 => D <= "11010111";	-- 0x05B2
		when 001459 => D <= "11010010";	-- 0x05B3
		when 001460 => D <= "11010010";	-- 0x05B4
		when 001461 => D <= "11010000";	-- 0x05B5
		when 001462 => D <= "11010000";	-- 0x05B6
		when 001463 => D <= "11010111";	-- 0x05B7
		when 001464 => D <= "00000000";	-- 0x05B8
		when 001465 => D <= "00000000";	-- 0x05B9
		when 001466 => D <= "11111100";	-- 0x05BA
		when 001467 => D <= "11111011";	-- 0x05BB
		when 001468 => D <= "11111001";	-- 0x05BC
		when 001469 => D <= "11111100";	-- 0x05BD
		when 001470 => D <= "00000000";	-- 0x05BE
		when 001471 => D <= "00000000";	-- 0x05BF
		when 001472 => D <= "00000000";	-- 0x05C0
		when 001473 => D <= "00000000";	-- 0x05C1
		when 001474 => D <= "11010101";	-- 0x05C2
		when 001475 => D <= "11010110";	-- 0x05C3
		when 001476 => D <= "11010110";	-- 0x05C4
		when 001477 => D <= "11010010";	-- 0x05C5
		when 001478 => D <= "11010010";	-- 0x05C6
		when 001479 => D <= "11010101";	-- 0x05C7
		when 001480 => D <= "00000000";	-- 0x05C8
		when 001481 => D <= "00000000";	-- 0x05C9
		when 001482 => D <= "11111000";	-- 0x05CA
		when 001483 => D <= "11111111";	-- 0x05CB
		when 001484 => D <= "11111011";	-- 0x05CC
		when 001485 => D <= "11111000";	-- 0x05CD
		when 001486 => D <= "00000000";	-- 0x05CE
		when 001487 => D <= "00000000";	-- 0x05CF
		when 001488 => D <= "00000000";	-- 0x05D0
		when 001489 => D <= "00000000";	-- 0x05D1
		when 001490 => D <= "11010001";	-- 0x05D2
		when 001491 => D <= "11010100";	-- 0x05D3
		when 001492 => D <= "11010100";	-- 0x05D4
		when 001493 => D <= "11010110";	-- 0x05D5
		when 001494 => D <= "11010110";	-- 0x05D6
		when 001495 => D <= "11010001";	-- 0x05D7
		when 001496 => D <= "00000000";	-- 0x05D8
		when 001497 => D <= "00000000";	-- 0x05D9
		when 001498 => D <= "11000101";	-- 0x05DA
		when 001499 => D <= "00000110";	-- 0x05DB
		when 001500 => D <= "00000100";	-- 0x05DC
		when 001501 => D <= "11001011";	-- 0x05DD
		when 001502 => D <= "00101100";	-- 0x05DE
		when 001503 => D <= "11001011";	-- 0x05DF
		when 001504 => D <= "00011101";	-- 0x05E0
		when 001505 => D <= "00000101";	-- 0x05E1
		when 001506 => D <= "11000010";	-- 0x05E2
		when 001507 => D <= "11011101";	-- 0x05E3
		when 001508 => D <= "00100101";	-- 0x05E4
		when 001509 => D <= "00111010";	-- 0x05E5
		when 001510 => D <= "01000100";	-- 0x05E6
		when 001511 => D <= "10000000";	-- 0x05E7
		when 001512 => D <= "11111110";	-- 0x05E8
		when 001513 => D <= "00000001";	-- 0x05E9
		when 001514 => D <= "11000010";	-- 0x05EA
		when 001515 => D <= "11110010";	-- 0x05EB
		when 001516 => D <= "00100101";	-- 0x05EC
		when 001517 => D <= "00000110";	-- 0x05ED
		when 001518 => D <= "00000101";	-- 0x05EE
		when 001519 => D <= "11000011";	-- 0x05EF
		when 001520 => D <= "11110100";	-- 0x05F0
		when 001521 => D <= "00100101";	-- 0x05F1
		when 001522 => D <= "00000110";	-- 0x05F2
		when 001523 => D <= "00000100";	-- 0x05F3
		when 001524 => D <= "11001011";	-- 0x05F4
		when 001525 => D <= "00101010";	-- 0x05F5
		when 001526 => D <= "11001011";	-- 0x05F6
		when 001527 => D <= "00011011";	-- 0x05F7
		when 001528 => D <= "00000101";	-- 0x05F8
		when 001529 => D <= "11000010";	-- 0x05F9
		when 001530 => D <= "11110100";	-- 0x05FA
		when 001531 => D <= "00100101";	-- 0x05FB
		when 001532 => D <= "11000001";	-- 0x05FC
		when 001533 => D <= "11001001";	-- 0x05FD
		when 001534 => D <= "11001101";	-- 0x05FE
		when 001535 => D <= "11100001";	-- 0x05FF
		when 001536 => D <= "00100110";	-- 0x0600
		when 001537 => D <= "11011000";	-- 0x0601
		when 001538 => D <= "11011101";	-- 0x0602
		when 001539 => D <= "01111110";	-- 0x0603
		when 001540 => D <= "00000000";	-- 0x0604
		when 001541 => D <= "11111110";	-- 0x0605
		when 001542 => D <= "00111100";	-- 0x0606
		when 001543 => D <= "11001010";	-- 0x0607
		when 001544 => D <= "00010100";	-- 0x0608
		when 001545 => D <= "00100110";	-- 0x0609
		when 001546 => D <= "11111110";	-- 0x060A
		when 001547 => D <= "00111110";	-- 0x060B
		when 001548 => D <= "11001010";	-- 0x060C
		when 001549 => D <= "00010100";	-- 0x060D
		when 001550 => D <= "00100110";	-- 0x060E
		when 001551 => D <= "11111110";	-- 0x060F
		when 001552 => D <= "00111101";	-- 0x0610
		when 001553 => D <= "11000010";	-- 0x0611
		when 001554 => D <= "11010101";	-- 0x0612
		when 001555 => D <= "00100110";	-- 0x0613
		when 001556 => D <= "11111110";	-- 0x0614
		when 001557 => D <= "00111101";	-- 0x0615
		when 001558 => D <= "11000010";	-- 0x0616
		when 001559 => D <= "00101111";	-- 0x0617
		when 001560 => D <= "00100110";	-- 0x0618
		when 001561 => D <= "11011101";	-- 0x0619
		when 001562 => D <= "00100011";	-- 0x061A
		when 001563 => D <= "11001101";	-- 0x061B
		when 001564 => D <= "11010111";	-- 0x061C
		when 001565 => D <= "00100110";	-- 0x061D
		when 001566 => D <= "01111100";	-- 0x061E
		when 001567 => D <= "10110101";	-- 0x061F
		when 001568 => D <= "11000010";	-- 0x0620
		when 001569 => D <= "00101001";	-- 0x0621
		when 001570 => D <= "00100110";	-- 0x0622
		when 001571 => D <= "00100001";	-- 0x0623
		when 001572 => D <= "11111111";	-- 0x0624
		when 001573 => D <= "11111111";	-- 0x0625
		when 001574 => D <= "11000011";	-- 0x0626
		when 001575 => D <= "00101100";	-- 0x0627
		when 001576 => D <= "00100110";	-- 0x0628
		when 001577 => D <= "00100001";	-- 0x0629
		when 001578 => D <= "00000000";	-- 0x062A
		when 001579 => D <= "00000000";	-- 0x062B
		when 001580 => D <= "11000011";	-- 0x062C
		when 001581 => D <= "11001111";	-- 0x062D
		when 001582 => D <= "00100110";	-- 0x062E
		when 001583 => D <= "11111110";	-- 0x062F
		when 001584 => D <= "00111100";	-- 0x0630
		when 001585 => D <= "11000010";	-- 0x0631
		when 001586 => D <= "10001100";	-- 0x0632
		when 001587 => D <= "00100110";	-- 0x0633
		when 001588 => D <= "11011101";	-- 0x0634
		when 001589 => D <= "01111110";	-- 0x0635
		when 001590 => D <= "00000001";	-- 0x0636
		when 001591 => D <= "11111110";	-- 0x0637
		when 001592 => D <= "00111101";	-- 0x0638
		when 001593 => D <= "11000010";	-- 0x0639
		when 001594 => D <= "01011111";	-- 0x063A
		when 001595 => D <= "00100110";	-- 0x063B
		when 001596 => D <= "11011101";	-- 0x063C
		when 001597 => D <= "00100011";	-- 0x063D
		when 001598 => D <= "11011101";	-- 0x063E
		when 001599 => D <= "00100011";	-- 0x063F
		when 001600 => D <= "11001101";	-- 0x0640
		when 001601 => D <= "11010111";	-- 0x0641
		when 001602 => D <= "00100110";	-- 0x0642
		when 001603 => D <= "11001011";	-- 0x0643
		when 001604 => D <= "01111100";	-- 0x0644
		when 001605 => D <= "11001010";	-- 0x0645
		when 001606 => D <= "01001110";	-- 0x0646
		when 001607 => D <= "00100110";	-- 0x0647
		when 001608 => D <= "00100001";	-- 0x0648
		when 001609 => D <= "11111111";	-- 0x0649
		when 001610 => D <= "11111111";	-- 0x064A
		when 001611 => D <= "11000011";	-- 0x064B
		when 001612 => D <= "01011100";	-- 0x064C
		when 001613 => D <= "00100110";	-- 0x064D
		when 001614 => D <= "01111100";	-- 0x064E
		when 001615 => D <= "10110101";	-- 0x064F
		when 001616 => D <= "11000010";	-- 0x0650
		when 001617 => D <= "01011001";	-- 0x0651
		when 001618 => D <= "00100110";	-- 0x0652
		when 001619 => D <= "00100001";	-- 0x0653
		when 001620 => D <= "11111111";	-- 0x0654
		when 001621 => D <= "11111111";	-- 0x0655
		when 001622 => D <= "11000011";	-- 0x0656
		when 001623 => D <= "01011100";	-- 0x0657
		when 001624 => D <= "00100110";	-- 0x0658
		when 001625 => D <= "00100001";	-- 0x0659
		when 001626 => D <= "00000000";	-- 0x065A
		when 001627 => D <= "00000000";	-- 0x065B
		when 001628 => D <= "11000011";	-- 0x065C
		when 001629 => D <= "10001001";	-- 0x065D
		when 001630 => D <= "00100110";	-- 0x065E
		when 001631 => D <= "11111110";	-- 0x065F
		when 001632 => D <= "00111110";	-- 0x0660
		when 001633 => D <= "11000010";	-- 0x0661
		when 001634 => D <= "01110110";	-- 0x0662
		when 001635 => D <= "00100110";	-- 0x0663
		when 001636 => D <= "11011101";	-- 0x0664
		when 001637 => D <= "00100011";	-- 0x0665
		when 001638 => D <= "11011101";	-- 0x0666
		when 001639 => D <= "00100011";	-- 0x0667
		when 001640 => D <= "11001101";	-- 0x0668
		when 001641 => D <= "11010111";	-- 0x0669
		when 001642 => D <= "00100110";	-- 0x066A
		when 001643 => D <= "01111100";	-- 0x066B
		when 001644 => D <= "10110101";	-- 0x066C
		when 001645 => D <= "11001010";	-- 0x066D
		when 001646 => D <= "01110011";	-- 0x066E
		when 001647 => D <= "00100110";	-- 0x066F
		when 001648 => D <= "00100001";	-- 0x0670
		when 001649 => D <= "11111111";	-- 0x0671
		when 001650 => D <= "11111111";	-- 0x0672
		when 001651 => D <= "11000011";	-- 0x0673
		when 001652 => D <= "10001001";	-- 0x0674
		when 001653 => D <= "00100110";	-- 0x0675
		when 001654 => D <= "11011101";	-- 0x0676
		when 001655 => D <= "00100011";	-- 0x0677
		when 001656 => D <= "11001101";	-- 0x0678
		when 001657 => D <= "11010111";	-- 0x0679
		when 001658 => D <= "00100110";	-- 0x067A
		when 001659 => D <= "11001011";	-- 0x067B
		when 001660 => D <= "01111100";	-- 0x067C
		when 001661 => D <= "11001010";	-- 0x067D
		when 001662 => D <= "10000110";	-- 0x067E
		when 001663 => D <= "00100110";	-- 0x067F
		when 001664 => D <= "00100001";	-- 0x0680
		when 001665 => D <= "11111111";	-- 0x0681
		when 001666 => D <= "11111111";	-- 0x0682
		when 001667 => D <= "11000011";	-- 0x0683
		when 001668 => D <= "10001001";	-- 0x0684
		when 001669 => D <= "00100110";	-- 0x0685
		when 001670 => D <= "00100001";	-- 0x0686
		when 001671 => D <= "00000000";	-- 0x0687
		when 001672 => D <= "00000000";	-- 0x0688
		when 001673 => D <= "11000011";	-- 0x0689
		when 001674 => D <= "11001111";	-- 0x068A
		when 001675 => D <= "00100110";	-- 0x068B
		when 001676 => D <= "11111110";	-- 0x068C
		when 001677 => D <= "00111110";	-- 0x068D
		when 001678 => D <= "11000010";	-- 0x068E
		when 001679 => D <= "11001111";	-- 0x068F
		when 001680 => D <= "00100110";	-- 0x0690
		when 001681 => D <= "11011101";	-- 0x0691
		when 001682 => D <= "01111110";	-- 0x0692
		when 001683 => D <= "00000001";	-- 0x0693
		when 001684 => D <= "11111110";	-- 0x0694
		when 001685 => D <= "00111101";	-- 0x0695
		when 001686 => D <= "11000010";	-- 0x0696
		when 001687 => D <= "10110001";	-- 0x0697
		when 001688 => D <= "00100110";	-- 0x0698
		when 001689 => D <= "11011101";	-- 0x0699
		when 001690 => D <= "00100011";	-- 0x069A
		when 001691 => D <= "11011101";	-- 0x069B
		when 001692 => D <= "00100011";	-- 0x069C
		when 001693 => D <= "11001101";	-- 0x069D
		when 001694 => D <= "11010111";	-- 0x069E
		when 001695 => D <= "00100110";	-- 0x069F
		when 001696 => D <= "11001011";	-- 0x06A0
		when 001697 => D <= "01111100";	-- 0x06A1
		when 001698 => D <= "11000010";	-- 0x06A2
		when 001699 => D <= "10101011";	-- 0x06A3
		when 001700 => D <= "00100110";	-- 0x06A4
		when 001701 => D <= "00100001";	-- 0x06A5
		when 001702 => D <= "11111111";	-- 0x06A6
		when 001703 => D <= "11111111";	-- 0x06A7
		when 001704 => D <= "11000011";	-- 0x06A8
		when 001705 => D <= "10101110";	-- 0x06A9
		when 001706 => D <= "00100110";	-- 0x06AA
		when 001707 => D <= "00100001";	-- 0x06AB
		when 001708 => D <= "00000000";	-- 0x06AC
		when 001709 => D <= "00000000";	-- 0x06AD
		when 001710 => D <= "11000011";	-- 0x06AE
		when 001711 => D <= "11001111";	-- 0x06AF
		when 001712 => D <= "00100110";	-- 0x06B0
		when 001713 => D <= "11011101";	-- 0x06B1
		when 001714 => D <= "00100011";	-- 0x06B2
		when 001715 => D <= "11001101";	-- 0x06B3
		when 001716 => D <= "11010111";	-- 0x06B4
		when 001717 => D <= "00100110";	-- 0x06B5
		when 001718 => D <= "11001011";	-- 0x06B6
		when 001719 => D <= "01111100";	-- 0x06B7
		when 001720 => D <= "11001010";	-- 0x06B8
		when 001721 => D <= "11000001";	-- 0x06B9
		when 001722 => D <= "00100110";	-- 0x06BA
		when 001723 => D <= "00100001";	-- 0x06BB
		when 001724 => D <= "00000000";	-- 0x06BC
		when 001725 => D <= "00000000";	-- 0x06BD
		when 001726 => D <= "11000011";	-- 0x06BE
		when 001727 => D <= "11001111";	-- 0x06BF
		when 001728 => D <= "00100110";	-- 0x06C0
		when 001729 => D <= "01111100";	-- 0x06C1
		when 001730 => D <= "10110101";	-- 0x06C2
		when 001731 => D <= "11000010";	-- 0x06C3
		when 001732 => D <= "11001100";	-- 0x06C4
		when 001733 => D <= "00100110";	-- 0x06C5
		when 001734 => D <= "00100001";	-- 0x06C6
		when 001735 => D <= "00000000";	-- 0x06C7
		when 001736 => D <= "00000000";	-- 0x06C8
		when 001737 => D <= "11000011";	-- 0x06C9
		when 001738 => D <= "11001111";	-- 0x06CA
		when 001739 => D <= "00100110";	-- 0x06CB
		when 001740 => D <= "00100001";	-- 0x06CC
		when 001741 => D <= "11111111";	-- 0x06CD
		when 001742 => D <= "11111111";	-- 0x06CE
		when 001743 => D <= "11011101";	-- 0x06CF
		when 001744 => D <= "01111110";	-- 0x06D0
		when 001745 => D <= "00000000";	-- 0x06D1
		when 001746 => D <= "11000011";	-- 0x06D2
		when 001747 => D <= "00000101";	-- 0x06D3
		when 001748 => D <= "00100110";	-- 0x06D4
		when 001749 => D <= "10101111";	-- 0x06D5
		when 001750 => D <= "11001001";	-- 0x06D6
		when 001751 => D <= "11100101";	-- 0x06D7
		when 001752 => D <= "11001101";	-- 0x06D8
		when 001753 => D <= "11100001";	-- 0x06D9
		when 001754 => D <= "00100110";	-- 0x06DA
		when 001755 => D <= "11010001";	-- 0x06DB
		when 001756 => D <= "11101011";	-- 0x06DC
		when 001757 => D <= "10101111";	-- 0x06DD
		when 001758 => D <= "11101101";	-- 0x06DE
		when 001759 => D <= "01010010";	-- 0x06DF
		when 001760 => D <= "11001001";	-- 0x06E0
		when 001761 => D <= "11001101";	-- 0x06E1
		when 001762 => D <= "00101111";	-- 0x06E2
		when 001763 => D <= "00100111";	-- 0x06E3
		when 001764 => D <= "11011000";	-- 0x06E4
		when 001765 => D <= "11011101";	-- 0x06E5
		when 001766 => D <= "01111110";	-- 0x06E6
		when 001767 => D <= "00000000";	-- 0x06E7
		when 001768 => D <= "11111110";	-- 0x06E8
		when 001769 => D <= "00101011";	-- 0x06E9
		when 001770 => D <= "11001010";	-- 0x06EA
		when 001771 => D <= "11110111";	-- 0x06EB
		when 001772 => D <= "00100110";	-- 0x06EC
		when 001773 => D <= "11111110";	-- 0x06ED
		when 001774 => D <= "00101101";	-- 0x06EE
		when 001775 => D <= "11001010";	-- 0x06EF
		when 001776 => D <= "11110111";	-- 0x06F0
		when 001777 => D <= "00100110";	-- 0x06F1
		when 001778 => D <= "11111110";	-- 0x06F2
		when 001779 => D <= "00100001";	-- 0x06F3
		when 001780 => D <= "11000010";	-- 0x06F4
		when 001781 => D <= "00101101";	-- 0x06F5
		when 001782 => D <= "00100111";	-- 0x06F6
		when 001783 => D <= "11011101";	-- 0x06F7
		when 001784 => D <= "00100011";	-- 0x06F8
		when 001785 => D <= "11111110";	-- 0x06F9
		when 001786 => D <= "00101011";	-- 0x06FA
		when 001787 => D <= "11000010";	-- 0x06FB
		when 001788 => D <= "00001000";	-- 0x06FC
		when 001789 => D <= "00100111";	-- 0x06FD
		when 001790 => D <= "11100101";	-- 0x06FE
		when 001791 => D <= "11001101";	-- 0x06FF
		when 001792 => D <= "00101111";	-- 0x0700
		when 001793 => D <= "00100111";	-- 0x0701
		when 001794 => D <= "11010001";	-- 0x0702
		when 001795 => D <= "11011000";	-- 0x0703
		when 001796 => D <= "00011001";	-- 0x0704
		when 001797 => D <= "11000011";	-- 0x0705
		when 001798 => D <= "00100111";	-- 0x0706
		when 001799 => D <= "00100111";	-- 0x0707
		when 001800 => D <= "11111110";	-- 0x0708
		when 001801 => D <= "00101101";	-- 0x0709
		when 001802 => D <= "11000010";	-- 0x070A
		when 001803 => D <= "00011010";	-- 0x070B
		when 001804 => D <= "00100111";	-- 0x070C
		when 001805 => D <= "11100101";	-- 0x070D
		when 001806 => D <= "11001101";	-- 0x070E
		when 001807 => D <= "00101111";	-- 0x070F
		when 001808 => D <= "00100111";	-- 0x0710
		when 001809 => D <= "11010001";	-- 0x0711
		when 001810 => D <= "11101011";	-- 0x0712
		when 001811 => D <= "11011000";	-- 0x0713
		when 001812 => D <= "10101111";	-- 0x0714
		when 001813 => D <= "11101101";	-- 0x0715
		when 001814 => D <= "01010010";	-- 0x0716
		when 001815 => D <= "11000011";	-- 0x0717
		when 001816 => D <= "00100111";	-- 0x0718
		when 001817 => D <= "00100111";	-- 0x0719
		when 001818 => D <= "11100101";	-- 0x071A
		when 001819 => D <= "11001101";	-- 0x071B
		when 001820 => D <= "00101111";	-- 0x071C
		when 001821 => D <= "00100111";	-- 0x071D
		when 001822 => D <= "11010001";	-- 0x071E
		when 001823 => D <= "11101011";	-- 0x071F
		when 001824 => D <= "11011000";	-- 0x0720
		when 001825 => D <= "01111101";	-- 0x0721
		when 001826 => D <= "10110011";	-- 0x0722
		when 001827 => D <= "01101111";	-- 0x0723
		when 001828 => D <= "01111100";	-- 0x0724
		when 001829 => D <= "10110100";	-- 0x0725
		when 001830 => D <= "01100111";	-- 0x0726
		when 001831 => D <= "11011101";	-- 0x0727
		when 001832 => D <= "01111110";	-- 0x0728
		when 001833 => D <= "00000000";	-- 0x0729
		when 001834 => D <= "11000011";	-- 0x072A
		when 001835 => D <= "11101000";	-- 0x072B
		when 001836 => D <= "00100110";	-- 0x072C
		when 001837 => D <= "10101111";	-- 0x072D
		when 001838 => D <= "11001001";	-- 0x072E
		when 001839 => D <= "11001101";	-- 0x072F
		when 001840 => D <= "11011101";	-- 0x0730
		when 001841 => D <= "00100111";	-- 0x0731
		when 001842 => D <= "11011000";	-- 0x0732
		when 001843 => D <= "11011101";	-- 0x0733
		when 001844 => D <= "01111110";	-- 0x0734
		when 001845 => D <= "00000000";	-- 0x0735
		when 001846 => D <= "11111110";	-- 0x0736
		when 001847 => D <= "00101010";	-- 0x0737
		when 001848 => D <= "11001010";	-- 0x0738
		when 001849 => D <= "01001010";	-- 0x0739
		when 001850 => D <= "00100111";	-- 0x073A
		when 001851 => D <= "11111110";	-- 0x073B
		when 001852 => D <= "00101111";	-- 0x073C
		when 001853 => D <= "11001010";	-- 0x073D
		when 001854 => D <= "01001010";	-- 0x073E
		when 001855 => D <= "00100111";	-- 0x073F
		when 001856 => D <= "11111110";	-- 0x0740
		when 001857 => D <= "01011100";	-- 0x0741
		when 001858 => D <= "11001010";	-- 0x0742
		when 001859 => D <= "01001010";	-- 0x0743
		when 001860 => D <= "00100111";	-- 0x0744
		when 001861 => D <= "11111110";	-- 0x0745
		when 001862 => D <= "00100110";	-- 0x0746
		when 001863 => D <= "11000010";	-- 0x0747
		when 001864 => D <= "11001010";	-- 0x0748
		when 001865 => D <= "00100111";	-- 0x0749
		when 001866 => D <= "11011101";	-- 0x074A
		when 001867 => D <= "00100011";	-- 0x074B
		when 001868 => D <= "11111110";	-- 0x074C
		when 001869 => D <= "00101010";	-- 0x074D
		when 001870 => D <= "11000010";	-- 0x074E
		when 001871 => D <= "01101011";	-- 0x074F
		when 001872 => D <= "00100111";	-- 0x0750
		when 001873 => D <= "11100101";	-- 0x0751
		when 001874 => D <= "11001101";	-- 0x0752
		when 001875 => D <= "11011101";	-- 0x0753
		when 001876 => D <= "00100111";	-- 0x0754
		when 001877 => D <= "11010001";	-- 0x0755
		when 001878 => D <= "11011000";	-- 0x0756
		when 001879 => D <= "11001101";	-- 0x0757
		when 001880 => D <= "10110110";	-- 0x0758
		when 001881 => D <= "00101001";	-- 0x0759
		when 001882 => D <= "11000101";	-- 0x075A
		when 001883 => D <= "11001101";	-- 0x075B
		when 001884 => D <= "11110010";	-- 0x075C
		when 001885 => D <= "00101001";	-- 0x075D
		when 001886 => D <= "11000001";	-- 0x075E
		when 001887 => D <= "01111000";	-- 0x075F
		when 001888 => D <= "11111110";	-- 0x0760
		when 001889 => D <= "00000001";	-- 0x0761
		when 001890 => D <= "11000010";	-- 0x0762
		when 001891 => D <= "01101000";	-- 0x0763
		when 001892 => D <= "00100111";	-- 0x0764
		when 001893 => D <= "11001101";	-- 0x0765
		when 001894 => D <= "11111010";	-- 0x0766
		when 001895 => D <= "00100010";	-- 0x0767
		when 001896 => D <= "11000011";	-- 0x0768
		when 001897 => D <= "11000100";	-- 0x0769
		when 001898 => D <= "00100111";	-- 0x076A
		when 001899 => D <= "11111110";	-- 0x076B
		when 001900 => D <= "00101111";	-- 0x076C
		when 001901 => D <= "11000010";	-- 0x076D
		when 001902 => D <= "10010001";	-- 0x076E
		when 001903 => D <= "00100111";	-- 0x076F
		when 001904 => D <= "11100101";	-- 0x0770
		when 001905 => D <= "11001101";	-- 0x0771
		when 001906 => D <= "11011101";	-- 0x0772
		when 001907 => D <= "00100111";	-- 0x0773
		when 001908 => D <= "11010001";	-- 0x0774
		when 001909 => D <= "11011000";	-- 0x0775
		when 001910 => D <= "11001101";	-- 0x0776
		when 001911 => D <= "10110110";	-- 0x0777
		when 001912 => D <= "00101001";	-- 0x0778
		when 001913 => D <= "11000101";	-- 0x0779
		when 001914 => D <= "01111011";	-- 0x077A
		when 001915 => D <= "10110010";	-- 0x077B
		when 001916 => D <= "11000010";	-- 0x077C
		when 001917 => D <= "10000001";	-- 0x077D
		when 001918 => D <= "00100111";	-- 0x077E
		when 001919 => D <= "00110111";	-- 0x077F
		when 001920 => D <= "11001001";	-- 0x0780
		when 001921 => D <= "11001101";	-- 0x0781
		when 001922 => D <= "11010000";	-- 0x0782
		when 001923 => D <= "00101001";	-- 0x0783
		when 001924 => D <= "11000001";	-- 0x0784
		when 001925 => D <= "01111000";	-- 0x0785
		when 001926 => D <= "11111110";	-- 0x0786
		when 001927 => D <= "00000001";	-- 0x0787
		when 001928 => D <= "11000010";	-- 0x0788
		when 001929 => D <= "10001110";	-- 0x0789
		when 001930 => D <= "00100111";	-- 0x078A
		when 001931 => D <= "11001101";	-- 0x078B
		when 001932 => D <= "11111010";	-- 0x078C
		when 001933 => D <= "00100010";	-- 0x078D
		when 001934 => D <= "11000011";	-- 0x078E
		when 001935 => D <= "11000100";	-- 0x078F
		when 001936 => D <= "00100111";	-- 0x0790
		when 001937 => D <= "11111110";	-- 0x0791
		when 001938 => D <= "01011100";	-- 0x0792
		when 001939 => D <= "11000010";	-- 0x0793
		when 001940 => D <= "10111000";	-- 0x0794
		when 001941 => D <= "00100111";	-- 0x0795
		when 001942 => D <= "11100101";	-- 0x0796
		when 001943 => D <= "11001101";	-- 0x0797
		when 001944 => D <= "11011101";	-- 0x0798
		when 001945 => D <= "00100111";	-- 0x0799
		when 001946 => D <= "11010001";	-- 0x079A
		when 001947 => D <= "11011000";	-- 0x079B
		when 001948 => D <= "11001101";	-- 0x079C
		when 001949 => D <= "10110110";	-- 0x079D
		when 001950 => D <= "00101001";	-- 0x079E
		when 001951 => D <= "11000101";	-- 0x079F
		when 001952 => D <= "01111011";	-- 0x07A0
		when 001953 => D <= "10110010";	-- 0x07A1
		when 001954 => D <= "11000010";	-- 0x07A2
		when 001955 => D <= "10100111";	-- 0x07A3
		when 001956 => D <= "00100111";	-- 0x07A4
		when 001957 => D <= "00110111";	-- 0x07A5
		when 001958 => D <= "11001001";	-- 0x07A6
		when 001959 => D <= "11001101";	-- 0x07A7
		when 001960 => D <= "11010000";	-- 0x07A8
		when 001961 => D <= "00101001";	-- 0x07A9
		when 001962 => D <= "11101011";	-- 0x07AA
		when 001963 => D <= "11000001";	-- 0x07AB
		when 001964 => D <= "01111000";	-- 0x07AC
		when 001965 => D <= "11111110";	-- 0x07AD
		when 001966 => D <= "00000001";	-- 0x07AE
		when 001967 => D <= "11000010";	-- 0x07AF
		when 001968 => D <= "10110101";	-- 0x07B0
		when 001969 => D <= "00100111";	-- 0x07B1
		when 001970 => D <= "11001101";	-- 0x07B2
		when 001971 => D <= "11111010";	-- 0x07B3
		when 001972 => D <= "00100010";	-- 0x07B4
		when 001973 => D <= "11000011";	-- 0x07B5
		when 001974 => D <= "11000100";	-- 0x07B6
		when 001975 => D <= "00100111";	-- 0x07B7
		when 001976 => D <= "11100101";	-- 0x07B8
		when 001977 => D <= "11001101";	-- 0x07B9
		when 001978 => D <= "11011101";	-- 0x07BA
		when 001979 => D <= "00100111";	-- 0x07BB
		when 001980 => D <= "11010001";	-- 0x07BC
		when 001981 => D <= "11011000";	-- 0x07BD
		when 001982 => D <= "01111101";	-- 0x07BE
		when 001983 => D <= "10100011";	-- 0x07BF
		when 001984 => D <= "01101111";	-- 0x07C0
		when 001985 => D <= "01111100";	-- 0x07C1
		when 001986 => D <= "10100010";	-- 0x07C2
		when 001987 => D <= "01100111";	-- 0x07C3
		when 001988 => D <= "11011101";	-- 0x07C4
		when 001989 => D <= "01111110";	-- 0x07C5
		when 001990 => D <= "00000000";	-- 0x07C6
		when 001991 => D <= "11000011";	-- 0x07C7
		when 001992 => D <= "00110110";	-- 0x07C8
		when 001993 => D <= "00100111";	-- 0x07C9
		when 001994 => D <= "10101111";	-- 0x07CA
		when 001995 => D <= "11001001";	-- 0x07CB
		when 001996 => D <= "11011101";	-- 0x07CC
		when 001997 => D <= "01111110";	-- 0x07CD
		when 001998 => D <= "00000000";	-- 0x07CE
		when 001999 => D <= "11111110";	-- 0x07CF
		when 002000 => D <= "00100000";	-- 0x07D0
		when 002001 => D <= "11000010";	-- 0x07D1
		when 002002 => D <= "11011100";	-- 0x07D2
		when 002003 => D <= "00100111";	-- 0x07D3
		when 002004 => D <= "11011101";	-- 0x07D4
		when 002005 => D <= "00100011";	-- 0x07D5
		when 002006 => D <= "11011101";	-- 0x07D6
		when 002007 => D <= "01111110";	-- 0x07D7
		when 002008 => D <= "00000000";	-- 0x07D8
		when 002009 => D <= "11000011";	-- 0x07D9
		when 002010 => D <= "11001111";	-- 0x07DA
		when 002011 => D <= "00100111";	-- 0x07DB
		when 002012 => D <= "11001001";	-- 0x07DC
		when 002013 => D <= "11011101";	-- 0x07DD
		when 002014 => D <= "01111110";	-- 0x07DE
		when 002015 => D <= "00000000";	-- 0x07DF
		when 002016 => D <= "11111110";	-- 0x07E0
		when 002017 => D <= "00101101";	-- 0x07E1
		when 002018 => D <= "11000010";	-- 0x07E2
		when 002019 => D <= "11110110";	-- 0x07E3
		when 002020 => D <= "00100111";	-- 0x07E4
		when 002021 => D <= "11011101";	-- 0x07E5
		when 002022 => D <= "00100011";	-- 0x07E6
		when 002023 => D <= "11001101";	-- 0x07E7
		when 002024 => D <= "11011101";	-- 0x07E8
		when 002025 => D <= "00100111";	-- 0x07E9
		when 002026 => D <= "11011000";	-- 0x07EA
		when 002027 => D <= "11101011";	-- 0x07EB
		when 002028 => D <= "00100001";	-- 0x07EC
		when 002029 => D <= "00000000";	-- 0x07ED
		when 002030 => D <= "00000000";	-- 0x07EE
		when 002031 => D <= "10101111";	-- 0x07EF
		when 002032 => D <= "11101101";	-- 0x07F0
		when 002033 => D <= "01010010";	-- 0x07F1
		when 002034 => D <= "10101111";	-- 0x07F2
		when 002035 => D <= "11000011";	-- 0x07F3
		when 002036 => D <= "01110011";	-- 0x07F4
		when 002037 => D <= "00101001";	-- 0x07F5
		when 002038 => D <= "11111110";	-- 0x07F6
		when 002039 => D <= "01111110";	-- 0x07F7
		when 002040 => D <= "11000010";	-- 0x07F8
		when 002041 => D <= "00001011";	-- 0x07F9
		when 002042 => D <= "00101000";	-- 0x07FA
		when 002043 => D <= "11011101";	-- 0x07FB
		when 002044 => D <= "00100011";	-- 0x07FC
		when 002045 => D <= "11001101";	-- 0x07FD
		when 002046 => D <= "11011101";	-- 0x07FE
		when 002047 => D <= "00100111";	-- 0x07FF
		when 002048 => D <= "11011000";	-- 0x0800
		when 002049 => D <= "01111100";	-- 0x0801
		when 002050 => D <= "00101111";	-- 0x0802
		when 002051 => D <= "01100111";	-- 0x0803
		when 002052 => D <= "01111101";	-- 0x0804
		when 002053 => D <= "00101111";	-- 0x0805
		when 002054 => D <= "01101111";	-- 0x0806
		when 002055 => D <= "10101111";	-- 0x0807
		when 002056 => D <= "11000011";	-- 0x0808
		when 002057 => D <= "01110011";	-- 0x0809
		when 002058 => D <= "00101001";	-- 0x080A
		when 002059 => D <= "11111110";	-- 0x080B
		when 002060 => D <= "00100010";	-- 0x080C
		when 002061 => D <= "11000010";	-- 0x080D
		when 002062 => D <= "00011100";	-- 0x080E
		when 002063 => D <= "00101000";	-- 0x080F
		when 002064 => D <= "11011101";	-- 0x0810
		when 002065 => D <= "00100011";	-- 0x0811
		when 002066 => D <= "11011101";	-- 0x0812
		when 002067 => D <= "01101110";	-- 0x0813
		when 002068 => D <= "00000000";	-- 0x0814
		when 002069 => D <= "00100110";	-- 0x0815
		when 002070 => D <= "00000000";	-- 0x0816
		when 002071 => D <= "11011101";	-- 0x0817
		when 002072 => D <= "00100011";	-- 0x0818
		when 002073 => D <= "11000011";	-- 0x0819
		when 002074 => D <= "01110011";	-- 0x081A
		when 002075 => D <= "00101001";	-- 0x081B
		when 002076 => D <= "11111110";	-- 0x081C
		when 002077 => D <= "00101000";	-- 0x081D
		when 002078 => D <= "11000010";	-- 0x081E
		when 002079 => D <= "00110101";	-- 0x081F
		when 002080 => D <= "00101000";	-- 0x0820
		when 002081 => D <= "11011101";	-- 0x0821
		when 002082 => D <= "00100011";	-- 0x0822
		when 002083 => D <= "11001101";	-- 0x0823
		when 002084 => D <= "11111110";	-- 0x0824
		when 002085 => D <= "00100101";	-- 0x0825
		when 002086 => D <= "11011101";	-- 0x0826
		when 002087 => D <= "01111110";	-- 0x0827
		when 002088 => D <= "00000000";	-- 0x0828
		when 002089 => D <= "11111110";	-- 0x0829
		when 002090 => D <= "00101001";	-- 0x082A
		when 002091 => D <= "11001010";	-- 0x082B
		when 002092 => D <= "00110000";	-- 0x082C
		when 002093 => D <= "00101000";	-- 0x082D
		when 002094 => D <= "00110111";	-- 0x082E
		when 002095 => D <= "11001001";	-- 0x082F
		when 002096 => D <= "11011101";	-- 0x0830
		when 002097 => D <= "00100011";	-- 0x0831
		when 002098 => D <= "11000011";	-- 0x0832
		when 002099 => D <= "01110011";	-- 0x0833
		when 002100 => D <= "00101001";	-- 0x0834
		when 002101 => D <= "11111110";	-- 0x0835
		when 002102 => D <= "00111010";	-- 0x0836
		when 002103 => D <= "11000010";	-- 0x0837
		when 002104 => D <= "01110000";	-- 0x0838
		when 002105 => D <= "00101001";	-- 0x0839
		when 002106 => D <= "11011101";	-- 0x083A
		when 002107 => D <= "00100011";	-- 0x083B
		when 002108 => D <= "11111101";	-- 0x083C
		when 002109 => D <= "00100001";	-- 0x083D
		when 002110 => D <= "01001111";	-- 0x083E
		when 002111 => D <= "10000011";	-- 0x083F
		when 002112 => D <= "11001101";	-- 0x0840
		when 002113 => D <= "00110101";	-- 0x0841
		when 002114 => D <= "00101010";	-- 0x0842
		when 002115 => D <= "11010010";	-- 0x0843
		when 002116 => D <= "01101101";	-- 0x0844
		when 002117 => D <= "00101001";	-- 0x0845
		when 002118 => D <= "11111101";	-- 0x0846
		when 002119 => D <= "00100001";	-- 0x0847
		when 002120 => D <= "01110100";	-- 0x0848
		when 002121 => D <= "00101001";	-- 0x0849
		when 002122 => D <= "11001101";	-- 0x084A
		when 002123 => D <= "00110101";	-- 0x084B
		when 002124 => D <= "00101010";	-- 0x084C
		when 002125 => D <= "11011010";	-- 0x084D
		when 002126 => D <= "01101101";	-- 0x084E
		when 002127 => D <= "00101001";	-- 0x084F
		when 002128 => D <= "01111101";	-- 0x0850
		when 002129 => D <= "11111110";	-- 0x0851
		when 002130 => D <= "00000001";	-- 0x0852
		when 002131 => D <= "11000010";	-- 0x0853
		when 002132 => D <= "01110010";	-- 0x0854
		when 002133 => D <= "00101000";	-- 0x0855
		when 002134 => D <= "11011101";	-- 0x0856
		when 002135 => D <= "01111110";	-- 0x0857
		when 002136 => D <= "00000000";	-- 0x0858
		when 002137 => D <= "11111110";	-- 0x0859
		when 002138 => D <= "00111111";	-- 0x085A
		when 002139 => D <= "11000010";	-- 0x085B
		when 002140 => D <= "01101000";	-- 0x085C
		when 002141 => D <= "00101000";	-- 0x085D
		when 002142 => D <= "11011101";	-- 0x085E
		when 002143 => D <= "00100011";	-- 0x085F
		when 002144 => D <= "11001101";	-- 0x0860
		when 002145 => D <= "00000011";	-- 0x0861
		when 002146 => D <= "00100000";	-- 0x0862
		when 002147 => D <= "01101111";	-- 0x0863
		when 002148 => D <= "01100101";	-- 0x0864
		when 002149 => D <= "11000011";	-- 0x0865
		when 002150 => D <= "01101110";	-- 0x0866
		when 002151 => D <= "00101000";	-- 0x0867
		when 002152 => D <= "11001101";	-- 0x0868
		when 002153 => D <= "00101001";	-- 0x0869
		when 002154 => D <= "00100000";	-- 0x086A
		when 002155 => D <= "01101111";	-- 0x086B
		when 002156 => D <= "00100110";	-- 0x086C
		when 002157 => D <= "00000000";	-- 0x086D
		when 002158 => D <= "10101111";	-- 0x086E
		when 002159 => D <= "11000011";	-- 0x086F
		when 002160 => D <= "01101101";	-- 0x0870
		when 002161 => D <= "00101001";	-- 0x0871
		when 002162 => D <= "11111110";	-- 0x0872
		when 002163 => D <= "00000010";	-- 0x0873
		when 002164 => D <= "11000010";	-- 0x0874
		when 002165 => D <= "10000010";	-- 0x0875
		when 002166 => D <= "00101000";	-- 0x0876
		when 002167 => D <= "11001101";	-- 0x0877
		when 002168 => D <= "00100010";	-- 0x0878
		when 002169 => D <= "00111100";	-- 0x0879
		when 002170 => D <= "01001101";	-- 0x087A
		when 002171 => D <= "11101101";	-- 0x087B
		when 002172 => D <= "01101000";	-- 0x087C
		when 002173 => D <= "00100110";	-- 0x087D
		when 002174 => D <= "00000000";	-- 0x087E
		when 002175 => D <= "11000011";	-- 0x087F
		when 002176 => D <= "01101101";	-- 0x0880
		when 002177 => D <= "00101001";	-- 0x0881
		when 002178 => D <= "11111110";	-- 0x0882
		when 002179 => D <= "00000011";	-- 0x0883
		when 002180 => D <= "11000010";	-- 0x0884
		when 002181 => D <= "11001111";	-- 0x0885
		when 002182 => D <= "00101000";	-- 0x0886
		when 002183 => D <= "00100001";	-- 0x0887
		when 002184 => D <= "00000000";	-- 0x0888
		when 002185 => D <= "00000000";	-- 0x0889
		when 002186 => D <= "00111010";	-- 0x088A
		when 002187 => D <= "01001000";	-- 0x088B
		when 002188 => D <= "10000000";	-- 0x088C
		when 002189 => D <= "11110101";	-- 0x088D
		when 002190 => D <= "11001101";	-- 0x088E
		when 002191 => D <= "00101001";	-- 0x088F
		when 002192 => D <= "00100000";	-- 0x0890
		when 002193 => D <= "11111110";	-- 0x0891
		when 002194 => D <= "00001000";	-- 0x0892
		when 002195 => D <= "11001010";	-- 0x0893
		when 002196 => D <= "10101111";	-- 0x0894
		when 002197 => D <= "00101000";	-- 0x0895
		when 002198 => D <= "11111110";	-- 0x0896
		when 002199 => D <= "00001001";	-- 0x0897
		when 002200 => D <= "11001010";	-- 0x0898
		when 002201 => D <= "10101111";	-- 0x0899
		when 002202 => D <= "00101000";	-- 0x089A
		when 002203 => D <= "11111110";	-- 0x089B
		when 002204 => D <= "01111111";	-- 0x089C
		when 002205 => D <= "11001010";	-- 0x089D
		when 002206 => D <= "10101111";	-- 0x089E
		when 002207 => D <= "00101000";	-- 0x089F
		when 002208 => D <= "11111110";	-- 0x08A0
		when 002209 => D <= "00000111";	-- 0x08A1
		when 002210 => D <= "11001010";	-- 0x08A2
		when 002211 => D <= "10101111";	-- 0x08A3
		when 002212 => D <= "00101000";	-- 0x08A4
		when 002213 => D <= "11111110";	-- 0x08A5
		when 002214 => D <= "10000000";	-- 0x08A6
		when 002215 => D <= "11010010";	-- 0x08A7
		when 002216 => D <= "10110011";	-- 0x08A8
		when 002217 => D <= "00101000";	-- 0x08A9
		when 002218 => D <= "11111110";	-- 0x08AA
		when 002219 => D <= "00100000";	-- 0x08AB
		when 002220 => D <= "11011010";	-- 0x08AC
		when 002221 => D <= "10110011";	-- 0x08AD
		when 002222 => D <= "00101000";	-- 0x08AE
		when 002223 => D <= "01001111";	-- 0x08AF
		when 002224 => D <= "11001101";	-- 0x08B0
		when 002225 => D <= "10110111";	-- 0x08B1
		when 002226 => D <= "00110000";	-- 0x08B2
		when 002227 => D <= "11111110";	-- 0x08B3
		when 002228 => D <= "00001101";	-- 0x08B4
		when 002229 => D <= "11000010";	-- 0x08B5
		when 002230 => D <= "10001110";	-- 0x08B6
		when 002231 => D <= "00101000";	-- 0x08B7
		when 002232 => D <= "11110001";	-- 0x08B8
		when 002233 => D <= "00110010";	-- 0x08B9
		when 002234 => D <= "01001000";	-- 0x08BA
		when 002235 => D <= "10000000";	-- 0x08BB
		when 002236 => D <= "11001101";	-- 0x08BC
		when 002237 => D <= "10111101";	-- 0x08BD
		when 002238 => D <= "00101100";	-- 0x08BE
		when 002239 => D <= "11011101";	-- 0x08BF
		when 002240 => D <= "11100101";	-- 0x08C0
		when 002241 => D <= "11100101";	-- 0x08C1
		when 002242 => D <= "11011101";	-- 0x08C2
		when 002243 => D <= "11100001";	-- 0x08C3
		when 002244 => D <= "11001101";	-- 0x08C4
		when 002245 => D <= "11001100";	-- 0x08C5
		when 002246 => D <= "00100111";	-- 0x08C6
		when 002247 => D <= "11001101";	-- 0x08C7
		when 002248 => D <= "11111110";	-- 0x08C8
		when 002249 => D <= "00100101";	-- 0x08C9
		when 002250 => D <= "11011101";	-- 0x08CA
		when 002251 => D <= "11100001";	-- 0x08CB
		when 002252 => D <= "11000011";	-- 0x08CC
		when 002253 => D <= "01101101";	-- 0x08CD
		when 002254 => D <= "00101001";	-- 0x08CE
		when 002255 => D <= "11111110";	-- 0x08CF
		when 002256 => D <= "00000100";	-- 0x08D0
		when 002257 => D <= "11000010";	-- 0x08D1
		when 002258 => D <= "11101010";	-- 0x08D2
		when 002259 => D <= "00101000";	-- 0x08D3
		when 002260 => D <= "11001101";	-- 0x08D4
		when 002261 => D <= "00100010";	-- 0x08D5
		when 002262 => D <= "00111100";	-- 0x08D6
		when 002263 => D <= "11011000";	-- 0x08D7
		when 002264 => D <= "11001101";	-- 0x08D8
		when 002265 => D <= "10100101";	-- 0x08D9
		when 002266 => D <= "00100010";	-- 0x08DA
		when 002267 => D <= "11001101";	-- 0x08DB
		when 002268 => D <= "01110001";	-- 0x08DC
		when 002269 => D <= "00100011";	-- 0x08DD
		when 002270 => D <= "01111000";	-- 0x08DE
		when 002271 => D <= "11111110";	-- 0x08DF
		when 002272 => D <= "00000001";	-- 0x08E0
		when 002273 => D <= "11000010";	-- 0x08E1
		when 002274 => D <= "11100111";	-- 0x08E2
		when 002275 => D <= "00101000";	-- 0x08E3
		when 002276 => D <= "11001101";	-- 0x08E4
		when 002277 => D <= "11111010";	-- 0x08E5
		when 002278 => D <= "00100010";	-- 0x08E6
		when 002279 => D <= "11000011";	-- 0x08E7
		when 002280 => D <= "01101101";	-- 0x08E8
		when 002281 => D <= "00101001";	-- 0x08E9
		when 002282 => D <= "11111110";	-- 0x08EA
		when 002283 => D <= "00000101";	-- 0x08EB
		when 002284 => D <= "11000010";	-- 0x08EC
		when 002285 => D <= "00000101";	-- 0x08ED
		when 002286 => D <= "00101001";	-- 0x08EE
		when 002287 => D <= "11001101";	-- 0x08EF
		when 002288 => D <= "00100010";	-- 0x08F0
		when 002289 => D <= "00111100";	-- 0x08F1
		when 002290 => D <= "11011000";	-- 0x08F2
		when 002291 => D <= "11001101";	-- 0x08F3
		when 002292 => D <= "10100101";	-- 0x08F4
		when 002293 => D <= "00100010";	-- 0x08F5
		when 002294 => D <= "11001101";	-- 0x08F6
		when 002295 => D <= "01100001";	-- 0x08F7
		when 002296 => D <= "00100011";	-- 0x08F8
		when 002297 => D <= "01111000";	-- 0x08F9
		when 002298 => D <= "11111110";	-- 0x08FA
		when 002299 => D <= "00000001";	-- 0x08FB
		when 002300 => D <= "11000010";	-- 0x08FC
		when 002301 => D <= "00000010";	-- 0x08FD
		when 002302 => D <= "00101001";	-- 0x08FE
		when 002303 => D <= "11001101";	-- 0x08FF
		when 002304 => D <= "11111010";	-- 0x0900
		when 002305 => D <= "00100010";	-- 0x0901
		when 002306 => D <= "11000011";	-- 0x0902
		when 002307 => D <= "01101101";	-- 0x0903
		when 002308 => D <= "00101001";	-- 0x0904
		when 002309 => D <= "11111110";	-- 0x0905
		when 002310 => D <= "00000110";	-- 0x0906
		when 002311 => D <= "11000010";	-- 0x0907
		when 002312 => D <= "00110101";	-- 0x0908
		when 002313 => D <= "00101001";	-- 0x0909
		when 002314 => D <= "11001101";	-- 0x090A
		when 002315 => D <= "00100010";	-- 0x090B
		when 002316 => D <= "00111100";	-- 0x090C
		when 002317 => D <= "11011000";	-- 0x090D
		when 002318 => D <= "11100101";	-- 0x090E
		when 002319 => D <= "11101101";	-- 0x090F
		when 002320 => D <= "01011111";	-- 0x0910
		when 002321 => D <= "01011111";	-- 0x0911
		when 002322 => D <= "00010110";	-- 0x0912
		when 002323 => D <= "00000000";	-- 0x0913
		when 002324 => D <= "00101010";	-- 0x0914
		when 002325 => D <= "00010100";	-- 0x0915
		when 002326 => D <= "10000000";	-- 0x0916
		when 002327 => D <= "00100011";	-- 0x0917
		when 002328 => D <= "01111100";	-- 0x0918
		when 002329 => D <= "11100110";	-- 0x0919
		when 002330 => D <= "00001111";	-- 0x091A
		when 002331 => D <= "01100111";	-- 0x091B
		when 002332 => D <= "00100010";	-- 0x091C
		when 002333 => D <= "00010100";	-- 0x091D
		when 002334 => D <= "10000000";	-- 0x091E
		when 002335 => D <= "00011001";	-- 0x091F
		when 002336 => D <= "01000110";	-- 0x0920
		when 002337 => D <= "11101101";	-- 0x0921
		when 002338 => D <= "01011111";	-- 0x0922
		when 002339 => D <= "10000000";	-- 0x0923
		when 002340 => D <= "01011111";	-- 0x0924
		when 002341 => D <= "00010110";	-- 0x0925
		when 002342 => D <= "00000000";	-- 0x0926
		when 002343 => D <= "11100001";	-- 0x0927
		when 002344 => D <= "11001101";	-- 0x0928
		when 002345 => D <= "11110010";	-- 0x0929
		when 002346 => D <= "00101001";	-- 0x092A
		when 002347 => D <= "00010001";	-- 0x092B
		when 002348 => D <= "00000000";	-- 0x092C
		when 002349 => D <= "00000001";	-- 0x092D
		when 002350 => D <= "11001101";	-- 0x092E
		when 002351 => D <= "11010000";	-- 0x092F
		when 002352 => D <= "00101001";	-- 0x0930
		when 002353 => D <= "10101111";	-- 0x0931
		when 002354 => D <= "11000011";	-- 0x0932
		when 002355 => D <= "01101101";	-- 0x0933
		when 002356 => D <= "00101001";	-- 0x0934
		when 002357 => D <= "11111110";	-- 0x0935
		when 002358 => D <= "00000111";	-- 0x0936
		when 002359 => D <= "11000010";	-- 0x0937
		when 002360 => D <= "01000100";	-- 0x0938
		when 002361 => D <= "00101001";	-- 0x0939
		when 002362 => D <= "00101010";	-- 0x093A
		when 002363 => D <= "00110111";	-- 0x093B
		when 002364 => D <= "10000000";	-- 0x093C
		when 002365 => D <= "11001101";	-- 0x093D
		when 002366 => D <= "11011010";	-- 0x093E
		when 002367 => D <= "00100101";	-- 0x093F
		when 002368 => D <= "10101111";	-- 0x0940
		when 002369 => D <= "11000011";	-- 0x0941
		when 002370 => D <= "01101101";	-- 0x0942
		when 002371 => D <= "00101001";	-- 0x0943
		when 002372 => D <= "11111110";	-- 0x0944
		when 002373 => D <= "00001000";	-- 0x0945
		when 002374 => D <= "11000010";	-- 0x0946
		when 002375 => D <= "01010011";	-- 0x0947
		when 002376 => D <= "00101001";	-- 0x0948
		when 002377 => D <= "00101010";	-- 0x0949
		when 002378 => D <= "00111001";	-- 0x094A
		when 002379 => D <= "10000000";	-- 0x094B
		when 002380 => D <= "11001101";	-- 0x094C
		when 002381 => D <= "11011010";	-- 0x094D
		when 002382 => D <= "00100101";	-- 0x094E
		when 002383 => D <= "10101111";	-- 0x094F
		when 002384 => D <= "11000011";	-- 0x0950
		when 002385 => D <= "01101101";	-- 0x0951
		when 002386 => D <= "00101001";	-- 0x0952
		when 002387 => D <= "11111110";	-- 0x0953
		when 002388 => D <= "00001001";	-- 0x0954
		when 002389 => D <= "11000010";	-- 0x0955
		when 002390 => D <= "01011111";	-- 0x0956
		when 002391 => D <= "00101001";	-- 0x0957
		when 002392 => D <= "00101010";	-- 0x0958
		when 002393 => D <= "00111011";	-- 0x0959
		when 002394 => D <= "10000000";	-- 0x095A
		when 002395 => D <= "10101111";	-- 0x095B
		when 002396 => D <= "11000011";	-- 0x095C
		when 002397 => D <= "01101101";	-- 0x095D
		when 002398 => D <= "00101001";	-- 0x095E
		when 002399 => D <= "11111110";	-- 0x095F
		when 002400 => D <= "10100000";	-- 0x0960
		when 002401 => D <= "11000010";	-- 0x0961
		when 002402 => D <= "01101101";	-- 0x0962
		when 002403 => D <= "00101001";	-- 0x0963
		when 002404 => D <= "11001101";	-- 0x0964
		when 002405 => D <= "00100010";	-- 0x0965
		when 002406 => D <= "00111100";	-- 0x0966
		when 002407 => D <= "11011000";	-- 0x0967
		when 002408 => D <= "01111110";	-- 0x0968
		when 002409 => D <= "00100110";	-- 0x0969
		when 002410 => D <= "00000000";	-- 0x096A
		when 002411 => D <= "01101111";	-- 0x096B
		when 002412 => D <= "10101111";	-- 0x096C
		when 002413 => D <= "11000011";	-- 0x096D
		when 002414 => D <= "01110011";	-- 0x096E
		when 002415 => D <= "00101001";	-- 0x096F
		when 002416 => D <= "11001101";	-- 0x0970
		when 002417 => D <= "11100001";	-- 0x0971
		when 002418 => D <= "00101011";	-- 0x0972
		when 002419 => D <= "11001001";	-- 0x0973
		when 002420 => D <= "01010100";	-- 0x0974
		when 002421 => D <= "01000001";	-- 0x0975
		when 002422 => D <= "01010011";	-- 0x0976
		when 002423 => D <= "01010100";	-- 0x0977
		when 002424 => D <= "11000101";	-- 0x0978
		when 002425 => D <= "00000001";	-- 0x0979
		when 002426 => D <= "00000000";	-- 0x097A
		when 002427 => D <= "00000000";	-- 0x097B
		when 002428 => D <= "01010000";	-- 0x097C
		when 002429 => D <= "01001111";	-- 0x097D
		when 002430 => D <= "01010010";	-- 0x097E
		when 002431 => D <= "11010100";	-- 0x097F
		when 002432 => D <= "00000010";	-- 0x0980
		when 002433 => D <= "00000000";	-- 0x0981
		when 002434 => D <= "00000000";	-- 0x0982
		when 002435 => D <= "01011010";	-- 0x0983
		when 002436 => D <= "01000001";	-- 0x0984
		when 002437 => D <= "01001000";	-- 0x0985
		when 002438 => D <= "11001100";	-- 0x0986
		when 002439 => D <= "00000011";	-- 0x0987
		when 002440 => D <= "00000000";	-- 0x0988
		when 002441 => D <= "00000000";	-- 0x0989
		when 002442 => D <= "01010011";	-- 0x098A
		when 002443 => D <= "01001001";	-- 0x098B
		when 002444 => D <= "11001110";	-- 0x098C
		when 002445 => D <= "00000100";	-- 0x098D
		when 002446 => D <= "00000000";	-- 0x098E
		when 002447 => D <= "00000000";	-- 0x098F
		when 002448 => D <= "01000011";	-- 0x0990
		when 002449 => D <= "01001111";	-- 0x0991
		when 002450 => D <= "11010011";	-- 0x0992
		when 002451 => D <= "00000101";	-- 0x0993
		when 002452 => D <= "00000000";	-- 0x0994
		when 002453 => D <= "00000000";	-- 0x0995
		when 002454 => D <= "01011010";	-- 0x0996
		when 002455 => D <= "11011010";	-- 0x0997
		when 002456 => D <= "00000110";	-- 0x0998
		when 002457 => D <= "00000000";	-- 0x0999
		when 002458 => D <= "00000000";	-- 0x099A
		when 002459 => D <= "01011000";	-- 0x099B
		when 002460 => D <= "01001011";	-- 0x099C
		when 002461 => D <= "11001111";	-- 0x099D
		when 002462 => D <= "00000111";	-- 0x099E
		when 002463 => D <= "00000000";	-- 0x099F
		when 002464 => D <= "00000000";	-- 0x09A0
		when 002465 => D <= "01011001";	-- 0x09A1
		when 002466 => D <= "01001011";	-- 0x09A2
		when 002467 => D <= "11001111";	-- 0x09A3
		when 002468 => D <= "00001000";	-- 0x09A4
		when 002469 => D <= "00000000";	-- 0x09A5
		when 002470 => D <= "00000000";	-- 0x09A6
		when 002471 => D <= "01001011";	-- 0x09A7
		when 002472 => D <= "01010101";	-- 0x09A8
		when 002473 => D <= "01010010";	-- 0x09A9
		when 002474 => D <= "11010011";	-- 0x09AA
		when 002475 => D <= "00001001";	-- 0x09AB
		when 002476 => D <= "00000000";	-- 0x09AC
		when 002477 => D <= "00000000";	-- 0x09AD
		when 002478 => D <= "01001101";	-- 0x09AE
		when 002479 => D <= "01000101";	-- 0x09AF
		when 002480 => D <= "11001101";	-- 0x09B0
		when 002481 => D <= "10100000";	-- 0x09B1
		when 002482 => D <= "00000000";	-- 0x09B2
		when 002483 => D <= "00000000";	-- 0x09B3
		when 002484 => D <= "00000000";	-- 0x09B4
		when 002485 => D <= "00000000";	-- 0x09B5
		when 002486 => D <= "00000110";	-- 0x09B6
		when 002487 => D <= "00000000";	-- 0x09B7
		when 002488 => D <= "11001011";	-- 0x09B8
		when 002489 => D <= "01111100";	-- 0x09B9
		when 002490 => D <= "11001010";	-- 0x09BA
		when 002491 => D <= "11000010";	-- 0x09BB
		when 002492 => D <= "00101001";	-- 0x09BC
		when 002493 => D <= "11001011";	-- 0x09BD
		when 002494 => D <= "11000000";	-- 0x09BE
		when 002495 => D <= "11001101";	-- 0x09BF
		when 002496 => D <= "11111010";	-- 0x09C0
		when 002497 => D <= "00100010";	-- 0x09C1
		when 002498 => D <= "11101011";	-- 0x09C2
		when 002499 => D <= "11001011";	-- 0x09C3
		when 002500 => D <= "01111100";	-- 0x09C4
		when 002501 => D <= "11001010";	-- 0x09C5
		when 002502 => D <= "11001111";	-- 0x09C6
		when 002503 => D <= "00101001";	-- 0x09C7
		when 002504 => D <= "01111000";	-- 0x09C8
		when 002505 => D <= "11101110";	-- 0x09C9
		when 002506 => D <= "00000001";	-- 0x09CA
		when 002507 => D <= "01000111";	-- 0x09CB
		when 002508 => D <= "11001101";	-- 0x09CC
		when 002509 => D <= "11111010";	-- 0x09CD
		when 002510 => D <= "00100010";	-- 0x09CE
		when 002511 => D <= "11001001";	-- 0x09CF
		when 002512 => D <= "00111110";	-- 0x09D0
		when 002513 => D <= "00010000";	-- 0x09D1
		when 002514 => D <= "11010101";	-- 0x09D2
		when 002515 => D <= "11000001";	-- 0x09D3
		when 002516 => D <= "00010001";	-- 0x09D4
		when 002517 => D <= "00000000";	-- 0x09D5
		when 002518 => D <= "00000000";	-- 0x09D6
		when 002519 => D <= "11101011";	-- 0x09D7
		when 002520 => D <= "11110101";	-- 0x09D8
		when 002521 => D <= "11001011";	-- 0x09D9
		when 002522 => D <= "00100011";	-- 0x09DA
		when 002523 => D <= "11001011";	-- 0x09DB
		when 002524 => D <= "00010010";	-- 0x09DC
		when 002525 => D <= "11001011";	-- 0x09DD
		when 002526 => D <= "00010101";	-- 0x09DE
		when 002527 => D <= "11001011";	-- 0x09DF
		when 002528 => D <= "00010100";	-- 0x09E0
		when 002529 => D <= "11001011";	-- 0x09E1
		when 002530 => D <= "11000011";	-- 0x09E2
		when 002531 => D <= "10101111";	-- 0x09E3
		when 002532 => D <= "11101101";	-- 0x09E4
		when 002533 => D <= "01000010";	-- 0x09E5
		when 002534 => D <= "11010010";	-- 0x09E6
		when 002535 => D <= "11101100";	-- 0x09E7
		when 002536 => D <= "00101001";	-- 0x09E8
		when 002537 => D <= "00001001";	-- 0x09E9
		when 002538 => D <= "11001011";	-- 0x09EA
		when 002539 => D <= "10000011";	-- 0x09EB
		when 002540 => D <= "11110001";	-- 0x09EC
		when 002541 => D <= "00111101";	-- 0x09ED
		when 002542 => D <= "00100000";	-- 0x09EE
		when 002543 => D <= "11101000";	-- 0x09EF
		when 002544 => D <= "11101011";	-- 0x09F0
		when 002545 => D <= "11001001";	-- 0x09F1
		when 002546 => D <= "00111110";	-- 0x09F2
		when 002547 => D <= "00010000";	-- 0x09F3
		when 002548 => D <= "11010101";	-- 0x09F4
		when 002549 => D <= "11000001";	-- 0x09F5
		when 002550 => D <= "00010001";	-- 0x09F6
		when 002551 => D <= "00000000";	-- 0x09F7
		when 002552 => D <= "00000000";	-- 0x09F8
		when 002553 => D <= "11101011";	-- 0x09F9
		when 002554 => D <= "11110101";	-- 0x09FA
		when 002555 => D <= "11001011";	-- 0x09FB
		when 002556 => D <= "01000011";	-- 0x09FC
		when 002557 => D <= "11001010";	-- 0x09FD
		when 002558 => D <= "00000001";	-- 0x09FE
		when 002559 => D <= "00101010";	-- 0x09FF
		when 002560 => D <= "00001001";	-- 0x0A00
		when 002561 => D <= "11001011";	-- 0x0A01
		when 002562 => D <= "00101100";	-- 0x0A02
		when 002563 => D <= "11001011";	-- 0x0A03
		when 002564 => D <= "00011101";	-- 0x0A04
		when 002565 => D <= "11001011";	-- 0x0A05
		when 002566 => D <= "00011010";	-- 0x0A06
		when 002567 => D <= "11001011";	-- 0x0A07
		when 002568 => D <= "00011011";	-- 0x0A08
		when 002569 => D <= "11110001";	-- 0x0A09
		when 002570 => D <= "00111101";	-- 0x0A0A
		when 002571 => D <= "00100000";	-- 0x0A0B
		when 002572 => D <= "11101101";	-- 0x0A0C
		when 002573 => D <= "11101011";	-- 0x0A0D
		when 002574 => D <= "11001001";	-- 0x0A0E
		when 002575 => D <= "11001011";	-- 0x0A0F
		when 002576 => D <= "01111100";	-- 0x0A10
		when 002577 => D <= "11001010";	-- 0x0A11
		when 002578 => D <= "00011100";	-- 0x0A12
		when 002579 => D <= "00101010";	-- 0x0A13
		when 002580 => D <= "00001110";	-- 0x0A14
		when 002581 => D <= "00101101";	-- 0x0A15
		when 002582 => D <= "11001101";	-- 0x0A16
		when 002583 => D <= "10110111";	-- 0x0A17
		when 002584 => D <= "00110000";	-- 0x0A18
		when 002585 => D <= "11001101";	-- 0x0A19
		when 002586 => D <= "11111010";	-- 0x0A1A
		when 002587 => D <= "00100010";	-- 0x0A1B
		when 002588 => D <= "10101111";	-- 0x0A1C
		when 002589 => D <= "11110101";	-- 0x0A1D
		when 002590 => D <= "00010001";	-- 0x0A1E
		when 002591 => D <= "00001010";	-- 0x0A1F
		when 002592 => D <= "00000000";	-- 0x0A20
		when 002593 => D <= "11001101";	-- 0x0A21
		when 002594 => D <= "11010000";	-- 0x0A22
		when 002595 => D <= "00101001";	-- 0x0A23
		when 002596 => D <= "01111011";	-- 0x0A24
		when 002597 => D <= "11110110";	-- 0x0A25
		when 002598 => D <= "00110000";	-- 0x0A26
		when 002599 => D <= "11110101";	-- 0x0A27
		when 002600 => D <= "01111100";	-- 0x0A28
		when 002601 => D <= "10110101";	-- 0x0A29
		when 002602 => D <= "00100000";	-- 0x0A2A
		when 002603 => D <= "11110010";	-- 0x0A2B
		when 002604 => D <= "11110001";	-- 0x0A2C
		when 002605 => D <= "10110111";	-- 0x0A2D
		when 002606 => D <= "11001000";	-- 0x0A2E
		when 002607 => D <= "01001111";	-- 0x0A2F
		when 002608 => D <= "11001101";	-- 0x0A30
		when 002609 => D <= "10110111";	-- 0x0A31
		when 002610 => D <= "00110000";	-- 0x0A32
		when 002611 => D <= "00011000";	-- 0x0A33
		when 002612 => D <= "11110111";	-- 0x0A34
		when 002613 => D <= "11011101";	-- 0x0A35
		when 002614 => D <= "01111110";	-- 0x0A36
		when 002615 => D <= "00000000";	-- 0x0A37
		when 002616 => D <= "11001011";	-- 0x0A38
		when 002617 => D <= "10111111";	-- 0x0A39
		when 002618 => D <= "11001101";	-- 0x0A3A
		when 002619 => D <= "10111100";	-- 0x0A3B
		when 002620 => D <= "00101010";	-- 0x0A3C
		when 002621 => D <= "11011000";	-- 0x0A3D
		when 002622 => D <= "11100101";	-- 0x0A3E
		when 002623 => D <= "00100001";	-- 0x0A3F
		when 002624 => D <= "10111011";	-- 0x0A40
		when 002625 => D <= "00101010";	-- 0x0A41
		when 002626 => D <= "11100011";	-- 0x0A42
		when 002627 => D <= "11111101";	-- 0x0A43
		when 002628 => D <= "01111110";	-- 0x0A44
		when 002629 => D <= "00000000";	-- 0x0A45
		when 002630 => D <= "10110111";	-- 0x0A46
		when 002631 => D <= "11000010";	-- 0x0A47
		when 002632 => D <= "01001100";	-- 0x0A48
		when 002633 => D <= "00101010";	-- 0x0A49
		when 002634 => D <= "00110111";	-- 0x0A4A
		when 002635 => D <= "11001001";	-- 0x0A4B
		when 002636 => D <= "11111101";	-- 0x0A4C
		when 002637 => D <= "00100010";	-- 0x0A4D
		when 002638 => D <= "11101000";	-- 0x0A4E
		when 002639 => D <= "10000010";	-- 0x0A4F
		when 002640 => D <= "11011101";	-- 0x0A50
		when 002641 => D <= "00100010";	-- 0x0A51
		when 002642 => D <= "11101010";	-- 0x0A52
		when 002643 => D <= "10000010";	-- 0x0A53
		when 002644 => D <= "11111101";	-- 0x0A54
		when 002645 => D <= "01000110";	-- 0x0A55
		when 002646 => D <= "00000000";	-- 0x0A56
		when 002647 => D <= "11001011";	-- 0x0A57
		when 002648 => D <= "10111000";	-- 0x0A58
		when 002649 => D <= "11011101";	-- 0x0A59
		when 002650 => D <= "01111110";	-- 0x0A5A
		when 002651 => D <= "00000000";	-- 0x0A5B
		when 002652 => D <= "11001011";	-- 0x0A5C
		when 002653 => D <= "10111111";	-- 0x0A5D
		when 002654 => D <= "11001101";	-- 0x0A5E
		when 002655 => D <= "11010010";	-- 0x0A5F
		when 002656 => D <= "00101011";	-- 0x0A60
		when 002657 => D <= "10111000";	-- 0x0A61
		when 002658 => D <= "11000010";	-- 0x0A62
		when 002659 => D <= "10010100";	-- 0x0A63
		when 002660 => D <= "00101010";	-- 0x0A64
		when 002661 => D <= "11011101";	-- 0x0A65
		when 002662 => D <= "00100011";	-- 0x0A66
		when 002663 => D <= "11111101";	-- 0x0A67
		when 002664 => D <= "11001011";	-- 0x0A68
		when 002665 => D <= "00000000";	-- 0x0A69
		when 002666 => D <= "01111110";	-- 0x0A6A
		when 002667 => D <= "11001010";	-- 0x0A6B
		when 002668 => D <= "10001110";	-- 0x0A6C
		when 002669 => D <= "00101010";	-- 0x0A6D
		when 002670 => D <= "11011101";	-- 0x0A6E
		when 002671 => D <= "01111110";	-- 0x0A6F
		when 002672 => D <= "00000000";	-- 0x0A70
		when 002673 => D <= "11001011";	-- 0x0A71
		when 002674 => D <= "10111111";	-- 0x0A72
		when 002675 => D <= "11001101";	-- 0x0A73
		when 002676 => D <= "10111100";	-- 0x0A74
		when 002677 => D <= "00101010";	-- 0x0A75
		when 002678 => D <= "11010010";	-- 0x0A76
		when 002679 => D <= "10001010";	-- 0x0A77
		when 002680 => D <= "00101010";	-- 0x0A78
		when 002681 => D <= "11111101";	-- 0x0A79
		when 002682 => D <= "00100011";	-- 0x0A7A
		when 002683 => D <= "11111101";	-- 0x0A7B
		when 002684 => D <= "01101110";	-- 0x0A7C
		when 002685 => D <= "00000000";	-- 0x0A7D
		when 002686 => D <= "11111101";	-- 0x0A7E
		when 002687 => D <= "01100110";	-- 0x0A7F
		when 002688 => D <= "00000001";	-- 0x0A80
		when 002689 => D <= "11111101";	-- 0x0A81
		when 002690 => D <= "01111110";	-- 0x0A82
		when 002691 => D <= "00000010";	-- 0x0A83
		when 002692 => D <= "00110111";	-- 0x0A84
		when 002693 => D <= "00111111";	-- 0x0A85
		when 002694 => D <= "11001001";	-- 0x0A86
		when 002695 => D <= "11000011";	-- 0x0A87
		when 002696 => D <= "10001011";	-- 0x0A88
		when 002697 => D <= "00101010";	-- 0x0A89
		when 002698 => D <= "00110111";	-- 0x0A8A
		when 002699 => D <= "11000011";	-- 0x0A8B
		when 002700 => D <= "10010001";	-- 0x0A8C
		when 002701 => D <= "00101010";	-- 0x0A8D
		when 002702 => D <= "11111101";	-- 0x0A8E
		when 002703 => D <= "00100011";	-- 0x0A8F
		when 002704 => D <= "10101111";	-- 0x0A90
		when 002705 => D <= "11000011";	-- 0x0A91
		when 002706 => D <= "10010101";	-- 0x0A92
		when 002707 => D <= "00101010";	-- 0x0A93
		when 002708 => D <= "00110111";	-- 0x0A94
		when 002709 => D <= "11010010";	-- 0x0A95
		when 002710 => D <= "01010100";	-- 0x0A96
		when 002711 => D <= "00101010";	-- 0x0A97
		when 002712 => D <= "11011101";	-- 0x0A98
		when 002713 => D <= "00101010";	-- 0x0A99
		when 002714 => D <= "11101010";	-- 0x0A9A
		when 002715 => D <= "10000010";	-- 0x0A9B
		when 002716 => D <= "11111101";	-- 0x0A9C
		when 002717 => D <= "00101010";	-- 0x0A9D
		when 002718 => D <= "11101000";	-- 0x0A9E
		when 002719 => D <= "10000010";	-- 0x0A9F
		when 002720 => D <= "11111101";	-- 0x0AA0
		when 002721 => D <= "11001011";	-- 0x0AA1
		when 002722 => D <= "00000000";	-- 0x0AA2
		when 002723 => D <= "01111110";	-- 0x0AA3
		when 002724 => D <= "11000010";	-- 0x0AA4
		when 002725 => D <= "10110000";	-- 0x0AA5
		when 002726 => D <= "00101010";	-- 0x0AA6
		when 002727 => D <= "11111101";	-- 0x0AA7
		when 002728 => D <= "00100011";	-- 0x0AA8
		when 002729 => D <= "11111101";	-- 0x0AA9
		when 002730 => D <= "11001011";	-- 0x0AAA
		when 002731 => D <= "00000000";	-- 0x0AAB
		when 002732 => D <= "01111110";	-- 0x0AAC
		when 002733 => D <= "11000011";	-- 0x0AAD
		when 002734 => D <= "10100100";	-- 0x0AAE
		when 002735 => D <= "00101010";	-- 0x0AAF
		when 002736 => D <= "11111101";	-- 0x0AB0
		when 002737 => D <= "00100011";	-- 0x0AB1
		when 002738 => D <= "11111101";	-- 0x0AB2
		when 002739 => D <= "00100011";	-- 0x0AB3
		when 002740 => D <= "11111101";	-- 0x0AB4
		when 002741 => D <= "00100011";	-- 0x0AB5
		when 002742 => D <= "11111101";	-- 0x0AB6
		when 002743 => D <= "00100011";	-- 0x0AB7
		when 002744 => D <= "11000011";	-- 0x0AB8
		when 002745 => D <= "01000011";	-- 0x0AB9
		when 002746 => D <= "00101010";	-- 0x0ABA
		when 002747 => D <= "11001001";	-- 0x0ABB
		when 002748 => D <= "11111110";	-- 0x0ABC
		when 002749 => D <= "00111010";	-- 0x0ABD
		when 002750 => D <= "00110000";	-- 0x0ABE
		when 002751 => D <= "00000101";	-- 0x0ABF
		when 002752 => D <= "11111110";	-- 0x0AC0
		when 002753 => D <= "00110000";	-- 0x0AC1
		when 002754 => D <= "11010010";	-- 0x0AC2
		when 002755 => D <= "11011100";	-- 0x0AC3
		when 002756 => D <= "00101010";	-- 0x0AC4
		when 002757 => D <= "11111110";	-- 0x0AC5
		when 002758 => D <= "01011011";	-- 0x0AC6
		when 002759 => D <= "00110000";	-- 0x0AC7
		when 002760 => D <= "00000101";	-- 0x0AC8
		when 002761 => D <= "11111110";	-- 0x0AC9
		when 002762 => D <= "01000001";	-- 0x0ACA
		when 002763 => D <= "11010010";	-- 0x0ACB
		when 002764 => D <= "11011100";	-- 0x0ACC
		when 002765 => D <= "00101010";	-- 0x0ACD
		when 002766 => D <= "11111110";	-- 0x0ACE
		when 002767 => D <= "01111011";	-- 0x0ACF
		when 002768 => D <= "00110000";	-- 0x0AD0
		when 002769 => D <= "00000101";	-- 0x0AD1
		when 002770 => D <= "11111110";	-- 0x0AD2
		when 002771 => D <= "01100001";	-- 0x0AD3
		when 002772 => D <= "11010010";	-- 0x0AD4
		when 002773 => D <= "11011100";	-- 0x0AD5
		when 002774 => D <= "00101010";	-- 0x0AD6
		when 002775 => D <= "11111110";	-- 0x0AD7
		when 002776 => D <= "01011111";	-- 0x0AD8
		when 002777 => D <= "11000010";	-- 0x0AD9
		when 002778 => D <= "11100001";	-- 0x0ADA
		when 002779 => D <= "00101010";	-- 0x0ADB
		when 002780 => D <= "00110111";	-- 0x0ADC
		when 002781 => D <= "00111111";	-- 0x0ADD
		when 002782 => D <= "11000011";	-- 0x0ADE
		when 002783 => D <= "11100010";	-- 0x0ADF
		when 002784 => D <= "00101010";	-- 0x0AE0
		when 002785 => D <= "00110111";	-- 0x0AE1
		when 002786 => D <= "11001001";	-- 0x0AE2
		when 002787 => D <= "11111101";	-- 0x0AE3
		when 002788 => D <= "00100001";	-- 0x0AE4
		when 002789 => D <= "01001111";	-- 0x0AE5
		when 002790 => D <= "10000011";	-- 0x0AE6
		when 002791 => D <= "11001101";	-- 0x0AE7
		when 002792 => D <= "00110101";	-- 0x0AE8
		when 002793 => D <= "00101010";	-- 0x0AE9
		when 002794 => D <= "11011000";	-- 0x0AEA
		when 002795 => D <= "11100101";	-- 0x0AEB
		when 002796 => D <= "00101010";	-- 0x0AEC
		when 002797 => D <= "01000111";	-- 0x0AED
		when 002798 => D <= "10000011";	-- 0x0AEE
		when 002799 => D <= "00101011";	-- 0x0AEF
		when 002800 => D <= "00100010";	-- 0x0AF0
		when 002801 => D <= "01000111";	-- 0x0AF1
		when 002802 => D <= "10000011";	-- 0x0AF2
		when 002803 => D <= "00101010";	-- 0x0AF3
		when 002804 => D <= "11101000";	-- 0x0AF4
		when 002805 => D <= "10000010";	-- 0x0AF5
		when 002806 => D <= "00010001";	-- 0x0AF6
		when 002807 => D <= "00000000";	-- 0x0AF7
		when 002808 => D <= "00000000";	-- 0x0AF8
		when 002809 => D <= "11001011";	-- 0x0AF9
		when 002810 => D <= "01111110";	-- 0x0AFA
		when 002811 => D <= "11000010";	-- 0x0AFB
		when 002812 => D <= "00000101";	-- 0x0AFC
		when 002813 => D <= "00101011";	-- 0x0AFD
		when 002814 => D <= "00010011";	-- 0x0AFE
		when 002815 => D <= "00100011";	-- 0x0AFF
		when 002816 => D <= "11001011";	-- 0x0B00
		when 002817 => D <= "01111110";	-- 0x0B01
		when 002818 => D <= "11000011";	-- 0x0B02
		when 002819 => D <= "11111011";	-- 0x0B03
		when 002820 => D <= "00101010";	-- 0x0B04
		when 002821 => D <= "00100011";	-- 0x0B05
		when 002822 => D <= "00010011";	-- 0x0B06
		when 002823 => D <= "00100011";	-- 0x0B07
		when 002824 => D <= "00010011";	-- 0x0B08
		when 002825 => D <= "00100011";	-- 0x0B09
		when 002826 => D <= "00010011";	-- 0x0B0A
		when 002827 => D <= "00100011";	-- 0x0B0B
		when 002828 => D <= "00010011";	-- 0x0B0C
		when 002829 => D <= "11100101";	-- 0x0B0D
		when 002830 => D <= "00101010";	-- 0x0B0E
		when 002831 => D <= "01001001";	-- 0x0B0F
		when 002832 => D <= "10000011";	-- 0x0B10
		when 002833 => D <= "11000001";	-- 0x0B11
		when 002834 => D <= "11000101";	-- 0x0B12
		when 002835 => D <= "10101111";	-- 0x0B13
		when 002836 => D <= "11101101";	-- 0x0B14
		when 002837 => D <= "01000010";	-- 0x0B15
		when 002838 => D <= "01000100";	-- 0x0B16
		when 002839 => D <= "01001101";	-- 0x0B17
		when 002840 => D <= "00000011";	-- 0x0B18
		when 002841 => D <= "00101010";	-- 0x0B19
		when 002842 => D <= "01001001";	-- 0x0B1A
		when 002843 => D <= "10000011";	-- 0x0B1B
		when 002844 => D <= "10101111";	-- 0x0B1C
		when 002845 => D <= "11101101";	-- 0x0B1D
		when 002846 => D <= "01010010";	-- 0x0B1E
		when 002847 => D <= "00100010";	-- 0x0B1F
		when 002848 => D <= "01001001";	-- 0x0B20
		when 002849 => D <= "10000011";	-- 0x0B21
		when 002850 => D <= "11100001";	-- 0x0B22
		when 002851 => D <= "11101101";	-- 0x0B23
		when 002852 => D <= "01011011";	-- 0x0B24
		when 002853 => D <= "11101000";	-- 0x0B25
		when 002854 => D <= "10000010";	-- 0x0B26
		when 002855 => D <= "11101101";	-- 0x0B27
		when 002856 => D <= "10110000";	-- 0x0B28
		when 002857 => D <= "11100001";	-- 0x0B29
		when 002858 => D <= "11001001";	-- 0x0B2A
		when 002859 => D <= "00110010";	-- 0x0B2B
		when 002860 => D <= "11101110";	-- 0x0B2C
		when 002861 => D <= "10000010";	-- 0x0B2D
		when 002862 => D <= "11101011";	-- 0x0B2E
		when 002863 => D <= "11100101";	-- 0x0B2F
		when 002864 => D <= "00100001";	-- 0x0B30
		when 002865 => D <= "01101101";	-- 0x0B31
		when 002866 => D <= "00101011";	-- 0x0B32
		when 002867 => D <= "11100011";	-- 0x0B33
		when 002868 => D <= "11111101";	-- 0x0B34
		when 002869 => D <= "00100010";	-- 0x0B35
		when 002870 => D <= "11101100";	-- 0x0B36
		when 002871 => D <= "10000010";	-- 0x0B37
		when 002872 => D <= "11111101";	-- 0x0B38
		when 002873 => D <= "01111110";	-- 0x0B39
		when 002874 => D <= "00000000";	-- 0x0B3A
		when 002875 => D <= "10110111";	-- 0x0B3B
		when 002876 => D <= "11000010";	-- 0x0B3C
		when 002877 => D <= "01000001";	-- 0x0B3D
		when 002878 => D <= "00101011";	-- 0x0B3E
		when 002879 => D <= "00110111";	-- 0x0B3F
		when 002880 => D <= "11001001";	-- 0x0B40
		when 002881 => D <= "11111101";	-- 0x0B41
		when 002882 => D <= "11001011";	-- 0x0B42
		when 002883 => D <= "00000000";	-- 0x0B43
		when 002884 => D <= "01111110";	-- 0x0B44
		when 002885 => D <= "11111101";	-- 0x0B45
		when 002886 => D <= "00100011";	-- 0x0B46
		when 002887 => D <= "11001010";	-- 0x0B47
		when 002888 => D <= "01000001";	-- 0x0B48
		when 002889 => D <= "00101011";	-- 0x0B49
		when 002890 => D <= "11111101";	-- 0x0B4A
		when 002891 => D <= "01101110";	-- 0x0B4B
		when 002892 => D <= "00000000";	-- 0x0B4C
		when 002893 => D <= "11111101";	-- 0x0B4D
		when 002894 => D <= "00100011";	-- 0x0B4E
		when 002895 => D <= "11111101";	-- 0x0B4F
		when 002896 => D <= "01100110";	-- 0x0B50
		when 002897 => D <= "00000000";	-- 0x0B51
		when 002898 => D <= "11111101";	-- 0x0B52
		when 002899 => D <= "00100011";	-- 0x0B53
		when 002900 => D <= "10101111";	-- 0x0B54
		when 002901 => D <= "11101101";	-- 0x0B55
		when 002902 => D <= "01010010";	-- 0x0B56
		when 002903 => D <= "11111101";	-- 0x0B57
		when 002904 => D <= "01000110";	-- 0x0B58
		when 002905 => D <= "00000000";	-- 0x0B59
		when 002906 => D <= "11111101";	-- 0x0B5A
		when 002907 => D <= "00100011";	-- 0x0B5B
		when 002908 => D <= "01111101";	-- 0x0B5C
		when 002909 => D <= "10110100";	-- 0x0B5D
		when 002910 => D <= "11000010";	-- 0x0B5E
		when 002911 => D <= "01101010";	-- 0x0B5F
		when 002912 => D <= "00101011";	-- 0x0B60
		when 002913 => D <= "00111010";	-- 0x0B61
		when 002914 => D <= "11101110";	-- 0x0B62
		when 002915 => D <= "10000010";	-- 0x0B63
		when 002916 => D <= "10111000";	-- 0x0B64
		when 002917 => D <= "11000010";	-- 0x0B65
		when 002918 => D <= "01101010";	-- 0x0B66
		when 002919 => D <= "00101011";	-- 0x0B67
		when 002920 => D <= "10101111";	-- 0x0B68
		when 002921 => D <= "11001001";	-- 0x0B69
		when 002922 => D <= "11000011";	-- 0x0B6A
		when 002923 => D <= "00110100";	-- 0x0B6B
		when 002924 => D <= "00101011";	-- 0x0B6C
		when 002925 => D <= "11111101";	-- 0x0B6D
		when 002926 => D <= "00101010";	-- 0x0B6E
		when 002927 => D <= "11101100";	-- 0x0B6F
		when 002928 => D <= "10000010";	-- 0x0B70
		when 002929 => D <= "11001001";	-- 0x0B71
		when 002930 => D <= "00110010";	-- 0x0B72
		when 002931 => D <= "11101110";	-- 0x0B73
		when 002932 => D <= "10000010";	-- 0x0B74
		when 002933 => D <= "11111101";	-- 0x0B75
		when 002934 => D <= "00100001";	-- 0x0B76
		when 002935 => D <= "01001111";	-- 0x0B77
		when 002936 => D <= "10000011";	-- 0x0B78
		when 002937 => D <= "11100101";	-- 0x0B79
		when 002938 => D <= "11011101";	-- 0x0B7A
		when 002939 => D <= "11100101";	-- 0x0B7B
		when 002940 => D <= "11001101";	-- 0x0B7C
		when 002941 => D <= "00110101";	-- 0x0B7D
		when 002942 => D <= "00101010";	-- 0x0B7E
		when 002943 => D <= "11011010";	-- 0x0B7F
		when 002944 => D <= "10000110";	-- 0x0B80
		when 002945 => D <= "00101011";	-- 0x0B81
		when 002946 => D <= "11000001";	-- 0x0B82
		when 002947 => D <= "11000001";	-- 0x0B83
		when 002948 => D <= "00110111";	-- 0x0B84
		when 002949 => D <= "11001001";	-- 0x0B85
		when 002950 => D <= "11011101";	-- 0x0B86
		when 002951 => D <= "11100001";	-- 0x0B87
		when 002952 => D <= "11100001";	-- 0x0B88
		when 002953 => D <= "11011101";	-- 0x0B89
		when 002954 => D <= "01111110";	-- 0x0B8A
		when 002955 => D <= "00000000";	-- 0x0B8B
		when 002956 => D <= "11001101";	-- 0x0B8C
		when 002957 => D <= "10111100";	-- 0x0B8D
		when 002958 => D <= "00101010";	-- 0x0B8E
		when 002959 => D <= "11011000";	-- 0x0B8F
		when 002960 => D <= "11111101";	-- 0x0B90
		when 002961 => D <= "00101010";	-- 0x0B91
		when 002962 => D <= "01001001";	-- 0x0B92
		when 002963 => D <= "10000011";	-- 0x0B93
		when 002964 => D <= "11011101";	-- 0x0B94
		when 002965 => D <= "01111110";	-- 0x0B95
		when 002966 => D <= "00000000";	-- 0x0B96
		when 002967 => D <= "11001101";	-- 0x0B97
		when 002968 => D <= "11010010";	-- 0x0B98
		when 002969 => D <= "00101011";	-- 0x0B99
		when 002970 => D <= "11111101";	-- 0x0B9A
		when 002971 => D <= "01110111";	-- 0x0B9B
		when 002972 => D <= "00000000";	-- 0x0B9C
		when 002973 => D <= "11011101";	-- 0x0B9D
		when 002974 => D <= "00100011";	-- 0x0B9E
		when 002975 => D <= "11111101";	-- 0x0B9F
		when 002976 => D <= "00100011";	-- 0x0BA0
		when 002977 => D <= "11011101";	-- 0x0BA1
		when 002978 => D <= "01111110";	-- 0x0BA2
		when 002979 => D <= "00000000";	-- 0x0BA3
		when 002980 => D <= "11001101";	-- 0x0BA4
		when 002981 => D <= "10111100";	-- 0x0BA5
		when 002982 => D <= "00101010";	-- 0x0BA6
		when 002983 => D <= "11010010";	-- 0x0BA7
		when 002984 => D <= "10010100";	-- 0x0BA8
		when 002985 => D <= "00101011";	-- 0x0BA9
		when 002986 => D <= "11111101";	-- 0x0BAA
		when 002987 => D <= "00101011";	-- 0x0BAB
		when 002988 => D <= "11111101";	-- 0x0BAC
		when 002989 => D <= "11001011";	-- 0x0BAD
		when 002990 => D <= "00000000";	-- 0x0BAE
		when 002991 => D <= "11111110";	-- 0x0BAF
		when 002992 => D <= "11111101";	-- 0x0BB0
		when 002993 => D <= "01110101";	-- 0x0BB1
		when 002994 => D <= "00000001";	-- 0x0BB2
		when 002995 => D <= "11111101";	-- 0x0BB3
		when 002996 => D <= "01110100";	-- 0x0BB4
		when 002997 => D <= "00000010";	-- 0x0BB5
		when 002998 => D <= "00111010";	-- 0x0BB6
		when 002999 => D <= "11101110";	-- 0x0BB7
		when 003000 => D <= "10000010";	-- 0x0BB8
		when 003001 => D <= "11111101";	-- 0x0BB9
		when 003002 => D <= "01110111";	-- 0x0BBA
		when 003003 => D <= "00000011";	-- 0x0BBB
		when 003004 => D <= "11111101";	-- 0x0BBC
		when 003005 => D <= "00110110";	-- 0x0BBD
		when 003006 => D <= "00000100";	-- 0x0BBE
		when 003007 => D <= "00000000";	-- 0x0BBF
		when 003008 => D <= "00010001";	-- 0x0BC0
		when 003009 => D <= "00000100";	-- 0x0BC1
		when 003010 => D <= "00000000";	-- 0x0BC2
		when 003011 => D <= "11111101";	-- 0x0BC3
		when 003012 => D <= "00011001";	-- 0x0BC4
		when 003013 => D <= "11111101";	-- 0x0BC5
		when 003014 => D <= "00100010";	-- 0x0BC6
		when 003015 => D <= "01001001";	-- 0x0BC7
		when 003016 => D <= "10000011";	-- 0x0BC8
		when 003017 => D <= "00101010";	-- 0x0BC9
		when 003018 => D <= "01000111";	-- 0x0BCA
		when 003019 => D <= "10000011";	-- 0x0BCB
		when 003020 => D <= "00100011";	-- 0x0BCC
		when 003021 => D <= "00100010";	-- 0x0BCD
		when 003022 => D <= "01000111";	-- 0x0BCE
		when 003023 => D <= "10000011";	-- 0x0BCF
		when 003024 => D <= "10101111";	-- 0x0BD0
		when 003025 => D <= "11001001";	-- 0x0BD1
		when 003026 => D <= "11111110";	-- 0x0BD2
		when 003027 => D <= "01111011";	-- 0x0BD3
		when 003028 => D <= "11010010";	-- 0x0BD4
		when 003029 => D <= "11100000";	-- 0x0BD5
		when 003030 => D <= "00101011";	-- 0x0BD6
		when 003031 => D <= "11111110";	-- 0x0BD7
		when 003032 => D <= "01100001";	-- 0x0BD8
		when 003033 => D <= "11011010";	-- 0x0BD9
		when 003034 => D <= "11100000";	-- 0x0BDA
		when 003035 => D <= "00101011";	-- 0x0BDB
		when 003036 => D <= "11010110";	-- 0x0BDC
		when 003037 => D <= "01100001";	-- 0x0BDD
		when 003038 => D <= "11000110";	-- 0x0BDE
		when 003039 => D <= "01000001";	-- 0x0BDF
		when 003040 => D <= "11001001";	-- 0x0BE0
		when 003041 => D <= "11011101";	-- 0x0BE1
		when 003042 => D <= "01111110";	-- 0x0BE2
		when 003043 => D <= "00000000";	-- 0x0BE3
		when 003044 => D <= "11111110";	-- 0x0BE4
		when 003045 => D <= "00101101";	-- 0x0BE5
		when 003046 => D <= "11000010";	-- 0x0BE6
		when 003047 => D <= "11110000";	-- 0x0BE7
		when 003048 => D <= "00101011";	-- 0x0BE8
		when 003049 => D <= "11011101";	-- 0x0BE9
		when 003050 => D <= "00100011";	-- 0x0BEA
		when 003051 => D <= "00111110";	-- 0x0BEB
		when 003052 => D <= "00000001";	-- 0x0BEC
		when 003053 => D <= "11000011";	-- 0x0BED
		when 003054 => D <= "11111100";	-- 0x0BEE
		when 003055 => D <= "00101011";	-- 0x0BEF
		when 003056 => D <= "11111110";	-- 0x0BF0
		when 003057 => D <= "00101011";	-- 0x0BF1
		when 003058 => D <= "11000010";	-- 0x0BF2
		when 003059 => D <= "11111011";	-- 0x0BF3
		when 003060 => D <= "00101011";	-- 0x0BF4
		when 003061 => D <= "11011101";	-- 0x0BF5
		when 003062 => D <= "00100011";	-- 0x0BF6
		when 003063 => D <= "10101111";	-- 0x0BF7
		when 003064 => D <= "11000011";	-- 0x0BF8
		when 003065 => D <= "11111100";	-- 0x0BF9
		when 003066 => D <= "00101011";	-- 0x0BFA
		when 003067 => D <= "10101111";	-- 0x0BFB
		when 003068 => D <= "00110010";	-- 0x0BFC
		when 003069 => D <= "00100100";	-- 0x0BFD
		when 003070 => D <= "10000000";	-- 0x0BFE
		when 003071 => D <= "00100001";	-- 0x0BFF
		when 003072 => D <= "00000000";	-- 0x0C00
		when 003073 => D <= "00000000";	-- 0x0C01
		when 003074 => D <= "11011101";	-- 0x0C02
		when 003075 => D <= "01111110";	-- 0x0C03
		when 003076 => D <= "00000000";	-- 0x0C04
		when 003077 => D <= "11001101";	-- 0x0C05
		when 003078 => D <= "00110110";	-- 0x0C06
		when 003079 => D <= "00101100";	-- 0x0C07
		when 003080 => D <= "11011000";	-- 0x0C08
		when 003081 => D <= "11011010";	-- 0x0C09
		when 003082 => D <= "00100011";	-- 0x0C0A
		when 003083 => D <= "00101100";	-- 0x0C0B
		when 003084 => D <= "11011101";	-- 0x0C0C
		when 003085 => D <= "00100011";	-- 0x0C0D
		when 003086 => D <= "01010100";	-- 0x0C0E
		when 003087 => D <= "01011101";	-- 0x0C0F
		when 003088 => D <= "00101001";	-- 0x0C10
		when 003089 => D <= "00101001";	-- 0x0C11
		when 003090 => D <= "00011001";	-- 0x0C12
		when 003091 => D <= "00101001";	-- 0x0C13
		when 003092 => D <= "11010110";	-- 0x0C14
		when 003093 => D <= "00110000";	-- 0x0C15
		when 003094 => D <= "01001111";	-- 0x0C16
		when 003095 => D <= "00000110";	-- 0x0C17
		when 003096 => D <= "00000000";	-- 0x0C18
		when 003097 => D <= "00001001";	-- 0x0C19
		when 003098 => D <= "11011101";	-- 0x0C1A
		when 003099 => D <= "01111110";	-- 0x0C1B
		when 003100 => D <= "00000000";	-- 0x0C1C
		when 003101 => D <= "11001101";	-- 0x0C1D
		when 003102 => D <= "00110110";	-- 0x0C1E
		when 003103 => D <= "00101100";	-- 0x0C1F
		when 003104 => D <= "11000011";	-- 0x0C20
		when 003105 => D <= "00001001";	-- 0x0C21
		when 003106 => D <= "00101100";	-- 0x0C22
		when 003107 => D <= "10101111";	-- 0x0C23
		when 003108 => D <= "11110101";	-- 0x0C24
		when 003109 => D <= "00111010";	-- 0x0C25
		when 003110 => D <= "00100100";	-- 0x0C26
		when 003111 => D <= "10000000";	-- 0x0C27
		when 003112 => D <= "11111110";	-- 0x0C28
		when 003113 => D <= "00000001";	-- 0x0C29
		when 003114 => D <= "11000010";	-- 0x0C2A
		when 003115 => D <= "00110100";	-- 0x0C2B
		when 003116 => D <= "00101100";	-- 0x0C2C
		when 003117 => D <= "11101011";	-- 0x0C2D
		when 003118 => D <= "00100001";	-- 0x0C2E
		when 003119 => D <= "00000000";	-- 0x0C2F
		when 003120 => D <= "00000000";	-- 0x0C30
		when 003121 => D <= "10101111";	-- 0x0C31
		when 003122 => D <= "11101101";	-- 0x0C32
		when 003123 => D <= "01010010";	-- 0x0C33
		when 003124 => D <= "11110001";	-- 0x0C34
		when 003125 => D <= "11001001";	-- 0x0C35
		when 003126 => D <= "11111110";	-- 0x0C36
		when 003127 => D <= "00111010";	-- 0x0C37
		when 003128 => D <= "11010010";	-- 0x0C38
		when 003129 => D <= "01000101";	-- 0x0C39
		when 003130 => D <= "00101100";	-- 0x0C3A
		when 003131 => D <= "11111110";	-- 0x0C3B
		when 003132 => D <= "00110000";	-- 0x0C3C
		when 003133 => D <= "11011010";	-- 0x0C3D
		when 003134 => D <= "01000101";	-- 0x0C3E
		when 003135 => D <= "00101100";	-- 0x0C3F
		when 003136 => D <= "00110111";	-- 0x0C40
		when 003137 => D <= "00111111";	-- 0x0C41
		when 003138 => D <= "11000011";	-- 0x0C42
		when 003139 => D <= "01000110";	-- 0x0C43
		when 003140 => D <= "00101100";	-- 0x0C44
		when 003141 => D <= "00110111";	-- 0x0C45
		when 003142 => D <= "11001001";	-- 0x0C46
		when 003143 => D <= "11100101";	-- 0x0C47
		when 003144 => D <= "11001101";	-- 0x0C48
		when 003145 => D <= "00010001";	-- 0x0C49
		when 003146 => D <= "00100001";	-- 0x0C4A
		when 003147 => D <= "00111110";	-- 0x0C4B
		when 003148 => D <= "00000000";	-- 0x0C4C
		when 003149 => D <= "00110010";	-- 0x0C4D
		when 003150 => D <= "01000110";	-- 0x0C4E
		when 003151 => D <= "10000000";	-- 0x0C4F
		when 003152 => D <= "00110010";	-- 0x0C50
		when 003153 => D <= "01000101";	-- 0x0C51
		when 003154 => D <= "10000000";	-- 0x0C52
		when 003155 => D <= "11001101";	-- 0x0C53
		when 003156 => D <= "01011000";	-- 0x0C54
		when 003157 => D <= "00100001";	-- 0x0C55
		when 003158 => D <= "00111110";	-- 0x0C56
		when 003159 => D <= "00000001";	-- 0x0C57
		when 003160 => D <= "00110010";	-- 0x0C58
		when 003161 => D <= "01000100";	-- 0x0C59
		when 003162 => D <= "10000000";	-- 0x0C5A
		when 003163 => D <= "00110010";	-- 0x0C5B
		when 003164 => D <= "01000011";	-- 0x0C5C
		when 003165 => D <= "10000000";	-- 0x0C5D
		when 003166 => D <= "00100001";	-- 0x0C5E
		when 003167 => D <= "00000000";	-- 0x0C5F
		when 003168 => D <= "00000000";	-- 0x0C60
		when 003169 => D <= "00100010";	-- 0x0C61
		when 003170 => D <= "00111101";	-- 0x0C62
		when 003171 => D <= "10000000";	-- 0x0C63
		when 003172 => D <= "00100010";	-- 0x0C64
		when 003173 => D <= "00111111";	-- 0x0C65
		when 003174 => D <= "10000000";	-- 0x0C66
		when 003175 => D <= "00100010";	-- 0x0C67
		when 003176 => D <= "01000001";	-- 0x0C68
		when 003177 => D <= "10000000";	-- 0x0C69
		when 003178 => D <= "00100010";	-- 0x0C6A
		when 003179 => D <= "00110111";	-- 0x0C6B
		when 003180 => D <= "10000000";	-- 0x0C6C
		when 003181 => D <= "00100010";	-- 0x0C6D
		when 003182 => D <= "00111001";	-- 0x0C6E
		when 003183 => D <= "10000000";	-- 0x0C6F
		when 003184 => D <= "00100010";	-- 0x0C70
		when 003185 => D <= "00111011";	-- 0x0C71
		when 003186 => D <= "10000000";	-- 0x0C72
		when 003187 => D <= "00111110";	-- 0x0C73
		when 003188 => D <= "00000001";	-- 0x0C74
		when 003189 => D <= "00110010";	-- 0x0C75
		when 003190 => D <= "00110110";	-- 0x0C76
		when 003191 => D <= "10000000";	-- 0x0C77
		when 003192 => D <= "11100001";	-- 0x0C78
		when 003193 => D <= "11001001";	-- 0x0C79
		when 003194 => D <= "00100001";	-- 0x0C7A
		when 003195 => D <= "01001011";	-- 0x0C7B
		when 003196 => D <= "10000011";	-- 0x0C7C
		when 003197 => D <= "01111110";	-- 0x0C7D
		when 003198 => D <= "00101111";	-- 0x0C7E
		when 003199 => D <= "01110111";	-- 0x0C7F
		when 003200 => D <= "10111110";	-- 0x0C80
		when 003201 => D <= "00100000";	-- 0x0C81
		when 003202 => D <= "00001101";	-- 0x0C82
		when 003203 => D <= "00101111";	-- 0x0C83
		when 003204 => D <= "01110111";	-- 0x0C84
		when 003205 => D <= "10111110";	-- 0x0C85
		when 003206 => D <= "00100000";	-- 0x0C86
		when 003207 => D <= "00001000";	-- 0x0C87
		when 003208 => D <= "00100011";	-- 0x0C88
		when 003209 => D <= "01111100";	-- 0x0C89
		when 003210 => D <= "11111110";	-- 0x0C8A
		when 003211 => D <= "11111111";	-- 0x0C8B
		when 003212 => D <= "00101000";	-- 0x0C8C
		when 003213 => D <= "00000010";	-- 0x0C8D
		when 003214 => D <= "00011000";	-- 0x0C8E
		when 003215 => D <= "11101101";	-- 0x0C8F
		when 003216 => D <= "00101011";	-- 0x0C90
		when 003217 => D <= "01000100";	-- 0x0C91
		when 003218 => D <= "01111101";	-- 0x0C92
		when 003219 => D <= "11001001";	-- 0x0C93
		when 003220 => D <= "11100101";	-- 0x0C94
		when 003221 => D <= "11010101";	-- 0x0C95
		when 003222 => D <= "00111010";	-- 0x0C96
		when 003223 => D <= "01001000";	-- 0x0C97
		when 003224 => D <= "10000000";	-- 0x0C98
		when 003225 => D <= "01001111";	-- 0x0C99
		when 003226 => D <= "01101001";	-- 0x0C9A
		when 003227 => D <= "00000110";	-- 0x0C9B
		when 003228 => D <= "00000000";	-- 0x0C9C
		when 003229 => D <= "01100000";	-- 0x0C9D
		when 003230 => D <= "00101001";	-- 0x0C9E
		when 003231 => D <= "00001001";	-- 0x0C9F
		when 003232 => D <= "00101001";	-- 0x0CA0
		when 003233 => D <= "11100101";	-- 0x0CA1
		when 003234 => D <= "00111010";	-- 0x0CA2
		when 003235 => D <= "01001001";	-- 0x0CA3
		when 003236 => D <= "10000000";	-- 0x0CA4
		when 003237 => D <= "01001111";	-- 0x0CA5
		when 003238 => D <= "01101001";	-- 0x0CA6
		when 003239 => D <= "00000110";	-- 0x0CA7
		when 003240 => D <= "00000000";	-- 0x0CA8
		when 003241 => D <= "01100000";	-- 0x0CA9
		when 003242 => D <= "00101001";	-- 0x0CAA
		when 003243 => D <= "00101001";	-- 0x0CAB
		when 003244 => D <= "00001001";	-- 0x0CAC
		when 003245 => D <= "00101001";	-- 0x0CAD
		when 003246 => D <= "00010001";	-- 0x0CAE
		when 003247 => D <= "01000110";	-- 0x0CAF
		when 003248 => D <= "00000000";	-- 0x0CB0
		when 003249 => D <= "11101011";	-- 0x0CB1
		when 003250 => D <= "10101111";	-- 0x0CB2
		when 003251 => D <= "11101101";	-- 0x0CB3
		when 003252 => D <= "01010010";	-- 0x0CB4
		when 003253 => D <= "11101011";	-- 0x0CB5
		when 003254 => D <= "11100001";	-- 0x0CB6
		when 003255 => D <= "11001101";	-- 0x0CB7
		when 003256 => D <= "01111010";	-- 0x0CB8
		when 003257 => D <= "00100001";	-- 0x0CB9
		when 003258 => D <= "11010001";	-- 0x0CBA
		when 003259 => D <= "11100001";	-- 0x0CBB
		when 003260 => D <= "11001001";	-- 0x0CBC
		when 003261 => D <= "00111010";	-- 0x0CBD
		when 003262 => D <= "01001001";	-- 0x0CBE
		when 003263 => D <= "10000000";	-- 0x0CBF
		when 003264 => D <= "01000111";	-- 0x0CC0
		when 003265 => D <= "11001101";	-- 0x0CC1
		when 003266 => D <= "10000101";	-- 0x0CC2
		when 003267 => D <= "00101110";	-- 0x0CC3
		when 003268 => D <= "00111010";	-- 0x0CC4
		when 003269 => D <= "01001000";	-- 0x0CC5
		when 003270 => D <= "10000000";	-- 0x0CC6
		when 003271 => D <= "01011111";	-- 0x0CC7
		when 003272 => D <= "00010110";	-- 0x0CC8
		when 003273 => D <= "00000000";	-- 0x0CC9
		when 003274 => D <= "00011001";	-- 0x0CCA
		when 003275 => D <= "11001001";	-- 0x0CCB
		when 003276 => D <= "11001101";	-- 0x0CCC
		when 003277 => D <= "10111101";	-- 0x0CCD
		when 003278 => D <= "00101100";	-- 0x0CCE
		when 003279 => D <= "01001110";	-- 0x0CCF
		when 003280 => D <= "11000101";	-- 0x0CD0
		when 003281 => D <= "11001101";	-- 0x0CD1
		when 003282 => D <= "01000010";	-- 0x0CD2
		when 003283 => D <= "00100010";	-- 0x0CD3
		when 003284 => D <= "00111110";	-- 0x0CD4
		when 003285 => D <= "00000000";	-- 0x0CD5
		when 003286 => D <= "00110010";	-- 0x0CD6
		when 003287 => D <= "01000110";	-- 0x0CD7
		when 003288 => D <= "10000000";	-- 0x0CD8
		when 003289 => D <= "11001101";	-- 0x0CD9
		when 003290 => D <= "01011000";	-- 0x0CDA
		when 003291 => D <= "00100001";	-- 0x0CDB
		when 003292 => D <= "11001101";	-- 0x0CDC
		when 003293 => D <= "10010100";	-- 0x0CDD
		when 003294 => D <= "00101100";	-- 0x0CDE
		when 003295 => D <= "00111110";	-- 0x0CDF
		when 003296 => D <= "00001010";	-- 0x0CE0
		when 003297 => D <= "11001101";	-- 0x0CE1
		when 003298 => D <= "11110011";	-- 0x0CE2
		when 003299 => D <= "00100000";	-- 0x0CE3
		when 003300 => D <= "11001101";	-- 0x0CE4
		when 003301 => D <= "10010100";	-- 0x0CE5
		when 003302 => D <= "00101100";	-- 0x0CE6
		when 003303 => D <= "11001101";	-- 0x0CE7
		when 003304 => D <= "01000110";	-- 0x0CE8
		when 003305 => D <= "00100010";	-- 0x0CE9
		when 003306 => D <= "11000001";	-- 0x0CEA
		when 003307 => D <= "01111001";	-- 0x0CEB
		when 003308 => D <= "11001101";	-- 0x0CEC
		when 003309 => D <= "11110011";	-- 0x0CED
		when 003310 => D <= "00100000";	-- 0x0CEE
		when 003311 => D <= "11001001";	-- 0x0CEF
		when 003312 => D <= "11001101";	-- 0x0CF0
		when 003313 => D <= "10111101";	-- 0x0CF1
		when 003314 => D <= "00101100";	-- 0x0CF2
		when 003315 => D <= "01111110";	-- 0x0CF3
		when 003316 => D <= "11110101";	-- 0x0CF4
		when 003317 => D <= "10101111";	-- 0x0CF5
		when 003318 => D <= "00110010";	-- 0x0CF6
		when 003319 => D <= "01000101";	-- 0x0CF7
		when 003320 => D <= "10000000";	-- 0x0CF8
		when 003321 => D <= "00110010";	-- 0x0CF9
		when 003322 => D <= "01000110";	-- 0x0CFA
		when 003323 => D <= "10000000";	-- 0x0CFB
		when 003324 => D <= "11001101";	-- 0x0CFC
		when 003325 => D <= "01011000";	-- 0x0CFD
		when 003326 => D <= "00100001";	-- 0x0CFE
		when 003327 => D <= "11001101";	-- 0x0CFF
		when 003328 => D <= "10010100";	-- 0x0D00
		when 003329 => D <= "00101100";	-- 0x0D01
		when 003330 => D <= "11001101";	-- 0x0D02
		when 003331 => D <= "01000110";	-- 0x0D03
		when 003332 => D <= "00100010";	-- 0x0D04
		when 003333 => D <= "00111110";	-- 0x0D05
		when 003334 => D <= "00001010";	-- 0x0D06
		when 003335 => D <= "11001101";	-- 0x0D07
		when 003336 => D <= "11110011";	-- 0x0D08
		when 003337 => D <= "00100000";	-- 0x0D09
		when 003338 => D <= "11001101";	-- 0x0D0A
		when 003339 => D <= "10010100";	-- 0x0D0B
		when 003340 => D <= "00101100";	-- 0x0D0C
		when 003341 => D <= "11001101";	-- 0x0D0D
		when 003342 => D <= "01000010";	-- 0x0D0E
		when 003343 => D <= "00100010";	-- 0x0D0F
		when 003344 => D <= "11110001";	-- 0x0D10
		when 003345 => D <= "11001101";	-- 0x0D11
		when 003346 => D <= "11110011";	-- 0x0D12
		when 003347 => D <= "00100000";	-- 0x0D13
		when 003348 => D <= "11001001";	-- 0x0D14
		when 003349 => D <= "00111010";	-- 0x0D15
		when 003350 => D <= "01010010";	-- 0x0D16
		when 003351 => D <= "10000000";	-- 0x0D17
		when 003352 => D <= "11110101";	-- 0x0D18
		when 003353 => D <= "11011101";	-- 0x0D19
		when 003354 => D <= "00100001";	-- 0x0D1A
		when 003355 => D <= "01010010";	-- 0x0D1B
		when 003356 => D <= "10000000";	-- 0x0D1C
		when 003357 => D <= "00000110";	-- 0x0D1D
		when 003358 => D <= "00000111";	-- 0x0D1E
		when 003359 => D <= "11011101";	-- 0x0D1F
		when 003360 => D <= "01111110";	-- 0x0D20
		when 003361 => D <= "00000001";	-- 0x0D21
		when 003362 => D <= "11011101";	-- 0x0D22
		when 003363 => D <= "01110111";	-- 0x0D23
		when 003364 => D <= "00000000";	-- 0x0D24
		when 003365 => D <= "11011101";	-- 0x0D25
		when 003366 => D <= "00100011";	-- 0x0D26
		when 003367 => D <= "00000101";	-- 0x0D27
		when 003368 => D <= "11000010";	-- 0x0D28
		when 003369 => D <= "00011111";	-- 0x0D29
		when 003370 => D <= "00101101";	-- 0x0D2A
		when 003371 => D <= "11110001";	-- 0x0D2B
		when 003372 => D <= "11011101";	-- 0x0D2C
		when 003373 => D <= "01110111";	-- 0x0D2D
		when 003374 => D <= "00000000";	-- 0x0D2E
		when 003375 => D <= "11001001";	-- 0x0D2F
		when 003376 => D <= "10101111";	-- 0x0D30
		when 003377 => D <= "00110010";	-- 0x0D31
		when 003378 => D <= "01000101";	-- 0x0D32
		when 003379 => D <= "10000000";	-- 0x0D33
		when 003380 => D <= "00111100";	-- 0x0D34
		when 003381 => D <= "00110010";	-- 0x0D35
		when 003382 => D <= "01000110";	-- 0x0D36
		when 003383 => D <= "10000000";	-- 0x0D37
		when 003384 => D <= "11001101";	-- 0x0D38
		when 003385 => D <= "01011000";	-- 0x0D39
		when 003386 => D <= "00100001";	-- 0x0D3A
		when 003387 => D <= "11001101";	-- 0x0D3B
		when 003388 => D <= "01000110";	-- 0x0D3C
		when 003389 => D <= "00100010";	-- 0x0D3D
		when 003390 => D <= "00100001";	-- 0x0D3E
		when 003391 => D <= "00000000";	-- 0x0D3F
		when 003392 => D <= "00000000";	-- 0x0D40
		when 003393 => D <= "00010001";	-- 0x0D41
		when 003394 => D <= "01000110";	-- 0x0D42
		when 003395 => D <= "00000000";	-- 0x0D43
		when 003396 => D <= "11001101";	-- 0x0D44
		when 003397 => D <= "01111010";	-- 0x0D45
		when 003398 => D <= "00100001";	-- 0x0D46
		when 003399 => D <= "11001101";	-- 0x0D47
		when 003400 => D <= "11011101";	-- 0x0D48
		when 003401 => D <= "00101110";	-- 0x0D49
		when 003402 => D <= "11001101";	-- 0x0D4A
		when 003403 => D <= "01000010";	-- 0x0D4B
		when 003404 => D <= "00100010";	-- 0x0D4C
		when 003405 => D <= "00100001";	-- 0x0D4D
		when 003406 => D <= "00000000";	-- 0x0D4E
		when 003407 => D <= "00000000";	-- 0x0D4F
		when 003408 => D <= "00010001";	-- 0x0D50
		when 003409 => D <= "01000110";	-- 0x0D51
		when 003410 => D <= "00000000";	-- 0x0D52
		when 003411 => D <= "11001101";	-- 0x0D53
		when 003412 => D <= "01111010";	-- 0x0D54
		when 003413 => D <= "00100001";	-- 0x0D55
		when 003414 => D <= "11001101";	-- 0x0D56
		when 003415 => D <= "11001100";	-- 0x0D57
		when 003416 => D <= "00101110";	-- 0x0D58
		when 003417 => D <= "10101111";	-- 0x0D59
		when 003418 => D <= "00110010";	-- 0x0D5A
		when 003419 => D <= "01000110";	-- 0x0D5B
		when 003420 => D <= "10000000";	-- 0x0D5C
		when 003421 => D <= "00111100";	-- 0x0D5D
		when 003422 => D <= "00110010";	-- 0x0D5E
		when 003423 => D <= "01000101";	-- 0x0D5F
		when 003424 => D <= "10000000";	-- 0x0D60
		when 003425 => D <= "11001101";	-- 0x0D61
		when 003426 => D <= "01011000";	-- 0x0D62
		when 003427 => D <= "00100001";	-- 0x0D63
		when 003428 => D <= "11001101";	-- 0x0D64
		when 003429 => D <= "01000110";	-- 0x0D65
		when 003430 => D <= "00100010";	-- 0x0D66
		when 003431 => D <= "00100001";	-- 0x0D67
		when 003432 => D <= "00000000";	-- 0x0D68
		when 003433 => D <= "00000000";	-- 0x0D69
		when 003434 => D <= "00010001";	-- 0x0D6A
		when 003435 => D <= "01000110";	-- 0x0D6B
		when 003436 => D <= "00000000";	-- 0x0D6C
		when 003437 => D <= "11001101";	-- 0x0D6D
		when 003438 => D <= "01111010";	-- 0x0D6E
		when 003439 => D <= "00100001";	-- 0x0D6F
		when 003440 => D <= "11001101";	-- 0x0D70
		when 003441 => D <= "11011101";	-- 0x0D71
		when 003442 => D <= "00101110";	-- 0x0D72
		when 003443 => D <= "11001101";	-- 0x0D73
		when 003444 => D <= "01000010";	-- 0x0D74
		when 003445 => D <= "00100010";	-- 0x0D75
		when 003446 => D <= "00100001";	-- 0x0D76
		when 003447 => D <= "00000000";	-- 0x0D77
		when 003448 => D <= "00000000";	-- 0x0D78
		when 003449 => D <= "00010001";	-- 0x0D79
		when 003450 => D <= "01000110";	-- 0x0D7A
		when 003451 => D <= "00000000";	-- 0x0D7B
		when 003452 => D <= "11001101";	-- 0x0D7C
		when 003453 => D <= "01111010";	-- 0x0D7D
		when 003454 => D <= "00100001";	-- 0x0D7E
		when 003455 => D <= "11001101";	-- 0x0D7F
		when 003456 => D <= "11001100";	-- 0x0D80
		when 003457 => D <= "00101110";	-- 0x0D81
		when 003458 => D <= "11001101";	-- 0x0D82
		when 003459 => D <= "00010101";	-- 0x0D83
		when 003460 => D <= "00101101";	-- 0x0D84
		when 003461 => D <= "00000110";	-- 0x0D85
		when 003462 => D <= "00000111";	-- 0x0D86
		when 003463 => D <= "11001101";	-- 0x0D87
		when 003464 => D <= "10000101";	-- 0x0D88
		when 003465 => D <= "00101110";	-- 0x0D89
		when 003466 => D <= "10101111";	-- 0x0D8A
		when 003467 => D <= "00000010";	-- 0x0D8B
		when 003468 => D <= "01010100";	-- 0x0D8C
		when 003469 => D <= "01011101";	-- 0x0D8D
		when 003470 => D <= "00010011";	-- 0x0D8E
		when 003471 => D <= "00000001";	-- 0x0D8F
		when 003472 => D <= "01001111";	-- 0x0D90
		when 003473 => D <= "00000000";	-- 0x0D91
		when 003474 => D <= "00110110";	-- 0x0D92
		when 003475 => D <= "00100000";	-- 0x0D93
		when 003476 => D <= "11101101";	-- 0x0D94
		when 003477 => D <= "10110000";	-- 0x0D95
		when 003478 => D <= "11001001";	-- 0x0D96
		when 003479 => D <= "10101111";	-- 0x0D97
		when 003480 => D <= "00110010";	-- 0x0D98
		when 003481 => D <= "01000101";	-- 0x0D99
		when 003482 => D <= "10000000";	-- 0x0D9A
		when 003483 => D <= "00111110";	-- 0x0D9B
		when 003484 => D <= "00000001";	-- 0x0D9C
		when 003485 => D <= "00110010";	-- 0x0D9D
		when 003486 => D <= "01000110";	-- 0x0D9E
		when 003487 => D <= "10000000";	-- 0x0D9F
		when 003488 => D <= "11001001";	-- 0x0DA0
		when 003489 => D <= "00111110";	-- 0x0DA1
		when 003490 => D <= "00000001";	-- 0x0DA2
		when 003491 => D <= "00110010";	-- 0x0DA3
		when 003492 => D <= "01000101";	-- 0x0DA4
		when 003493 => D <= "10000000";	-- 0x0DA5
		when 003494 => D <= "10101111";	-- 0x0DA6
		when 003495 => D <= "00110010";	-- 0x0DA7
		when 003496 => D <= "01000110";	-- 0x0DA8
		when 003497 => D <= "10000000";	-- 0x0DA9
		when 003498 => D <= "11001001";	-- 0x0DAA
		when 003499 => D <= "11001101";	-- 0x0DAB
		when 003500 => D <= "10010111";	-- 0x0DAC
		when 003501 => D <= "00101101";	-- 0x0DAD
		when 003502 => D <= "11001101";	-- 0x0DAE
		when 003503 => D <= "01011000";	-- 0x0DAF
		when 003504 => D <= "00100001";	-- 0x0DB0
		when 003505 => D <= "11001101";	-- 0x0DB1
		when 003506 => D <= "10010100";	-- 0x0DB2
		when 003507 => D <= "00101100";	-- 0x0DB3
		when 003508 => D <= "11001101";	-- 0x0DB4
		when 003509 => D <= "01000110";	-- 0x0DB5
		when 003510 => D <= "00100010";	-- 0x0DB6
		when 003511 => D <= "11001101";	-- 0x0DB7
		when 003512 => D <= "10101100";	-- 0x0DB8
		when 003513 => D <= "00101110";	-- 0x0DB9
		when 003514 => D <= "11001101";	-- 0x0DBA
		when 003515 => D <= "10010100";	-- 0x0DBB
		when 003516 => D <= "00101100";	-- 0x0DBC
		when 003517 => D <= "11001101";	-- 0x0DBD
		when 003518 => D <= "01000010";	-- 0x0DBE
		when 003519 => D <= "00100010";	-- 0x0DBF
		when 003520 => D <= "00111110";	-- 0x0DC0
		when 003521 => D <= "00100000";	-- 0x0DC1
		when 003522 => D <= "11001101";	-- 0x0DC2
		when 003523 => D <= "11110011";	-- 0x0DC3
		when 003524 => D <= "00100000";	-- 0x0DC4
		when 003525 => D <= "00111010";	-- 0x0DC5
		when 003526 => D <= "01001000";	-- 0x0DC6
		when 003527 => D <= "10000000";	-- 0x0DC7
		when 003528 => D <= "11111110";	-- 0x0DC8
		when 003529 => D <= "01001111";	-- 0x0DC9
		when 003530 => D <= "11010010";	-- 0x0DCA
		when 003531 => D <= "11010000";	-- 0x0DCB
		when 003532 => D <= "00101101";	-- 0x0DCC
		when 003533 => D <= "11001101";	-- 0x0DCD
		when 003534 => D <= "10100101";	-- 0x0DCE
		when 003535 => D <= "00101110";	-- 0x0DCF
		when 003536 => D <= "11001101";	-- 0x0DD0
		when 003537 => D <= "10100001";	-- 0x0DD1
		when 003538 => D <= "00101101";	-- 0x0DD2
		when 003539 => D <= "11001101";	-- 0x0DD3
		when 003540 => D <= "01011000";	-- 0x0DD4
		when 003541 => D <= "00100001";	-- 0x0DD5
		when 003542 => D <= "11001101";	-- 0x0DD6
		when 003543 => D <= "10010100";	-- 0x0DD7
		when 003544 => D <= "00101100";	-- 0x0DD8
		when 003545 => D <= "11001101";	-- 0x0DD9
		when 003546 => D <= "01000110";	-- 0x0DDA
		when 003547 => D <= "00100010";	-- 0x0DDB
		when 003548 => D <= "11001101";	-- 0x0DDC
		when 003549 => D <= "10101100";	-- 0x0DDD
		when 003550 => D <= "00101110";	-- 0x0DDE
		when 003551 => D <= "11001101";	-- 0x0DDF
		when 003552 => D <= "10010100";	-- 0x0DE0
		when 003553 => D <= "00101100";	-- 0x0DE1
		when 003554 => D <= "11001101";	-- 0x0DE2
		when 003555 => D <= "01000010";	-- 0x0DE3
		when 003556 => D <= "00100010";	-- 0x0DE4
		when 003557 => D <= "00111110";	-- 0x0DE5
		when 003558 => D <= "00100000";	-- 0x0DE6
		when 003559 => D <= "11001101";	-- 0x0DE7
		when 003560 => D <= "11110011";	-- 0x0DE8
		when 003561 => D <= "00100000";	-- 0x0DE9
		when 003562 => D <= "00111010";	-- 0x0DEA
		when 003563 => D <= "01001000";	-- 0x0DEB
		when 003564 => D <= "10000000";	-- 0x0DEC
		when 003565 => D <= "11111110";	-- 0x0DED
		when 003566 => D <= "01001111";	-- 0x0DEE
		when 003567 => D <= "11010010";	-- 0x0DEF
		when 003568 => D <= "11110101";	-- 0x0DF0
		when 003569 => D <= "00101101";	-- 0x0DF1
		when 003570 => D <= "11001101";	-- 0x0DF2
		when 003571 => D <= "10100101";	-- 0x0DF3
		when 003572 => D <= "00101110";	-- 0x0DF4
		when 003573 => D <= "11001101";	-- 0x0DF5
		when 003574 => D <= "10111101";	-- 0x0DF6
		when 003575 => D <= "00101100";	-- 0x0DF7
		when 003576 => D <= "00001010";	-- 0x0DF8
		when 003577 => D <= "11111110";	-- 0x0DF9
		when 003578 => D <= "01010000";	-- 0x0DFA
		when 003579 => D <= "11010010";	-- 0x0DFB
		when 003580 => D <= "00000000";	-- 0x0DFC
		when 003581 => D <= "00101110";	-- 0x0DFD
		when 003582 => D <= "00111100";	-- 0x0DFE
		when 003583 => D <= "00000010";	-- 0x0DFF
		when 003584 => D <= "00111010";	-- 0x0E00
		when 003585 => D <= "01001000";	-- 0x0E01
		when 003586 => D <= "10000000";	-- 0x0E02
		when 003587 => D <= "01000111";	-- 0x0E03
		when 003588 => D <= "00001110";	-- 0x0E04
		when 003589 => D <= "00100000";	-- 0x0E05
		when 003590 => D <= "01111110";	-- 0x0E06
		when 003591 => D <= "01110001";	-- 0x0E07
		when 003592 => D <= "01001111";	-- 0x0E08
		when 003593 => D <= "00100011";	-- 0x0E09
		when 003594 => D <= "00000100";	-- 0x0E0A
		when 003595 => D <= "01111000";	-- 0x0E0B
		when 003596 => D <= "11111110";	-- 0x0E0C
		when 003597 => D <= "01010000";	-- 0x0E0D
		when 003598 => D <= "11000010";	-- 0x0E0E
		when 003599 => D <= "00000110";	-- 0x0E0F
		when 003600 => D <= "00101110";	-- 0x0E10
		when 003601 => D <= "11001001";	-- 0x0E11
		when 003602 => D <= "11001101";	-- 0x0E12
		when 003603 => D <= "10010111";	-- 0x0E13
		when 003604 => D <= "00101101";	-- 0x0E14
		when 003605 => D <= "11001101";	-- 0x0E15
		when 003606 => D <= "01011000";	-- 0x0E16
		when 003607 => D <= "00100001";	-- 0x0E17
		when 003608 => D <= "11001101";	-- 0x0E18
		when 003609 => D <= "10010100";	-- 0x0E19
		when 003610 => D <= "00101100";	-- 0x0E1A
		when 003611 => D <= "11001101";	-- 0x0E1B
		when 003612 => D <= "01000110";	-- 0x0E1C
		when 003613 => D <= "00100010";	-- 0x0E1D
		when 003614 => D <= "11001101";	-- 0x0E1E
		when 003615 => D <= "10101100";	-- 0x0E1F
		when 003616 => D <= "00101110";	-- 0x0E20
		when 003617 => D <= "11001101";	-- 0x0E21
		when 003618 => D <= "10010100";	-- 0x0E22
		when 003619 => D <= "00101100";	-- 0x0E23
		when 003620 => D <= "11001101";	-- 0x0E24
		when 003621 => D <= "01000010";	-- 0x0E25
		when 003622 => D <= "00100010";	-- 0x0E26
		when 003623 => D <= "00111010";	-- 0x0E27
		when 003624 => D <= "01001000";	-- 0x0E28
		when 003625 => D <= "10000000";	-- 0x0E29
		when 003626 => D <= "11110101";	-- 0x0E2A
		when 003627 => D <= "00111100";	-- 0x0E2B
		when 003628 => D <= "11111110";	-- 0x0E2C
		when 003629 => D <= "01010000";	-- 0x0E2D
		when 003630 => D <= "11010010";	-- 0x0E2E
		when 003631 => D <= "00110111";	-- 0x0E2F
		when 003632 => D <= "00101110";	-- 0x0E30
		when 003633 => D <= "00110010";	-- 0x0E31
		when 003634 => D <= "01001000";	-- 0x0E32
		when 003635 => D <= "10000000";	-- 0x0E33
		when 003636 => D <= "11001101";	-- 0x0E34
		when 003637 => D <= "10101100";	-- 0x0E35
		when 003638 => D <= "00101110";	-- 0x0E36
		when 003639 => D <= "11110001";	-- 0x0E37
		when 003640 => D <= "00110010";	-- 0x0E38
		when 003641 => D <= "01001000";	-- 0x0E39
		when 003642 => D <= "10000000";	-- 0x0E3A
		when 003643 => D <= "11001101";	-- 0x0E3B
		when 003644 => D <= "10100001";	-- 0x0E3C
		when 003645 => D <= "00101101";	-- 0x0E3D
		when 003646 => D <= "11001101";	-- 0x0E3E
		when 003647 => D <= "01011000";	-- 0x0E3F
		when 003648 => D <= "00100001";	-- 0x0E40
		when 003649 => D <= "11001101";	-- 0x0E41
		when 003650 => D <= "10010100";	-- 0x0E42
		when 003651 => D <= "00101100";	-- 0x0E43
		when 003652 => D <= "11001101";	-- 0x0E44
		when 003653 => D <= "01000110";	-- 0x0E45
		when 003654 => D <= "00100010";	-- 0x0E46
		when 003655 => D <= "11001101";	-- 0x0E47
		when 003656 => D <= "10101100";	-- 0x0E48
		when 003657 => D <= "00101110";	-- 0x0E49
		when 003658 => D <= "11001101";	-- 0x0E4A
		when 003659 => D <= "10010100";	-- 0x0E4B
		when 003660 => D <= "00101100";	-- 0x0E4C
		when 003661 => D <= "11001101";	-- 0x0E4D
		when 003662 => D <= "01000010";	-- 0x0E4E
		when 003663 => D <= "00100010";	-- 0x0E4F
		when 003664 => D <= "00111010";	-- 0x0E50
		when 003665 => D <= "01001000";	-- 0x0E51
		when 003666 => D <= "10000000";	-- 0x0E52
		when 003667 => D <= "11110101";	-- 0x0E53
		when 003668 => D <= "00111100";	-- 0x0E54
		when 003669 => D <= "11111110";	-- 0x0E55
		when 003670 => D <= "01010000";	-- 0x0E56
		when 003671 => D <= "11010010";	-- 0x0E57
		when 003672 => D <= "01100000";	-- 0x0E58
		when 003673 => D <= "00101110";	-- 0x0E59
		when 003674 => D <= "00110010";	-- 0x0E5A
		when 003675 => D <= "01001000";	-- 0x0E5B
		when 003676 => D <= "10000000";	-- 0x0E5C
		when 003677 => D <= "11001101";	-- 0x0E5D
		when 003678 => D <= "10101100";	-- 0x0E5E
		when 003679 => D <= "00101110";	-- 0x0E5F
		when 003680 => D <= "11110001";	-- 0x0E60
		when 003681 => D <= "00110010";	-- 0x0E61
		when 003682 => D <= "01001000";	-- 0x0E62
		when 003683 => D <= "10000000";	-- 0x0E63
		when 003684 => D <= "11001101";	-- 0x0E64
		when 003685 => D <= "10111101";	-- 0x0E65
		when 003686 => D <= "00101100";	-- 0x0E66
		when 003687 => D <= "00111010";	-- 0x0E67
		when 003688 => D <= "01001000";	-- 0x0E68
		when 003689 => D <= "10000000";	-- 0x0E69
		when 003690 => D <= "01000111";	-- 0x0E6A
		when 003691 => D <= "11100101";	-- 0x0E6B
		when 003692 => D <= "11011101";	-- 0x0E6C
		when 003693 => D <= "11100001";	-- 0x0E6D
		when 003694 => D <= "01111000";	-- 0x0E6E
		when 003695 => D <= "11111110";	-- 0x0E6F
		when 003696 => D <= "01001111";	-- 0x0E70
		when 003697 => D <= "11010010";	-- 0x0E71
		when 003698 => D <= "10000000";	-- 0x0E72
		when 003699 => D <= "00101110";	-- 0x0E73
		when 003700 => D <= "11011101";	-- 0x0E74
		when 003701 => D <= "01111110";	-- 0x0E75
		when 003702 => D <= "00000001";	-- 0x0E76
		when 003703 => D <= "11011101";	-- 0x0E77
		when 003704 => D <= "01110111";	-- 0x0E78
		when 003705 => D <= "00000000";	-- 0x0E79
		when 003706 => D <= "11011101";	-- 0x0E7A
		when 003707 => D <= "00100011";	-- 0x0E7B
		when 003708 => D <= "00000100";	-- 0x0E7C
		when 003709 => D <= "11000011";	-- 0x0E7D
		when 003710 => D <= "01101110";	-- 0x0E7E
		when 003711 => D <= "00101110";	-- 0x0E7F
		when 003712 => D <= "11011101";	-- 0x0E80
		when 003713 => D <= "00110110";	-- 0x0E81
		when 003714 => D <= "00000000";	-- 0x0E82
		when 003715 => D <= "00100000";	-- 0x0E83
		when 003716 => D <= "11001001";	-- 0x0E84
		when 003717 => D <= "11010101";	-- 0x0E85
		when 003718 => D <= "01011000";	-- 0x0E86
		when 003719 => D <= "00010110";	-- 0x0E87
		when 003720 => D <= "00000000";	-- 0x0E88
		when 003721 => D <= "00100001";	-- 0x0E89
		when 003722 => D <= "01010010";	-- 0x0E8A
		when 003723 => D <= "10000000";	-- 0x0E8B
		when 003724 => D <= "00011001";	-- 0x0E8C
		when 003725 => D <= "01011110";	-- 0x0E8D
		when 003726 => D <= "00100001";	-- 0x0E8E
		when 003727 => D <= "01001010";	-- 0x0E8F
		when 003728 => D <= "10000000";	-- 0x0E90
		when 003729 => D <= "00011001";	-- 0x0E91
		when 003730 => D <= "01000100";	-- 0x0E92
		when 003731 => D <= "01001101";	-- 0x0E93
		when 003732 => D <= "01100010";	-- 0x0E94
		when 003733 => D <= "01101011";	-- 0x0E95
		when 003734 => D <= "00101001";	-- 0x0E96
		when 003735 => D <= "00101001";	-- 0x0E97
		when 003736 => D <= "00101001";	-- 0x0E98
		when 003737 => D <= "00101001";	-- 0x0E99
		when 003738 => D <= "01010100";	-- 0x0E9A
		when 003739 => D <= "01011101";	-- 0x0E9B
		when 003740 => D <= "00101001";	-- 0x0E9C
		when 003741 => D <= "00101001";	-- 0x0E9D
		when 003742 => D <= "00011001";	-- 0x0E9E
		when 003743 => D <= "00010001";	-- 0x0E9F
		when 003744 => D <= "01011010";	-- 0x0EA0
		when 003745 => D <= "10000000";	-- 0x0EA1
		when 003746 => D <= "00011001";	-- 0x0EA2
		when 003747 => D <= "11010001";	-- 0x0EA3
		when 003748 => D <= "11001001";	-- 0x0EA4
		when 003749 => D <= "00111110";	-- 0x0EA5
		when 003750 => D <= "01001111";	-- 0x0EA6
		when 003751 => D <= "00110010";	-- 0x0EA7
		when 003752 => D <= "11011101";	-- 0x0EA8
		when 003753 => D <= "10000010";	-- 0x0EA9
		when 003754 => D <= "00011000";	-- 0x0EAA
		when 003755 => D <= "00000101";	-- 0x0EAB
		when 003756 => D <= "00111110";	-- 0x0EAC
		when 003757 => D <= "01010000";	-- 0x0EAD
		when 003758 => D <= "00110010";	-- 0x0EAE
		when 003759 => D <= "11011101";	-- 0x0EAF
		when 003760 => D <= "10000010";	-- 0x0EB0
		when 003761 => D <= "11001101";	-- 0x0EB1
		when 003762 => D <= "10111101";	-- 0x0EB2
		when 003763 => D <= "00101100";	-- 0x0EB3
		when 003764 => D <= "00111010";	-- 0x0EB4
		when 003765 => D <= "01001000";	-- 0x0EB5
		when 003766 => D <= "10000000";	-- 0x0EB6
		when 003767 => D <= "01001111";	-- 0x0EB7
		when 003768 => D <= "11011011";	-- 0x0EB8
		when 003769 => D <= "01110000";	-- 0x0EB9
		when 003770 => D <= "11100110";	-- 0x0EBA
		when 003771 => D <= "00000100";	-- 0x0EBB
		when 003772 => D <= "11001010";	-- 0x0EBC
		when 003773 => D <= "10111000";	-- 0x0EBD
		when 003774 => D <= "00101110";	-- 0x0EBE
		when 003775 => D <= "01111110";	-- 0x0EBF
		when 003776 => D <= "11010011";	-- 0x0EC0
		when 003777 => D <= "01110000";	-- 0x0EC1
		when 003778 => D <= "00100011";	-- 0x0EC2
		when 003779 => D <= "00001100";	-- 0x0EC3
		when 003780 => D <= "00111010";	-- 0x0EC4
		when 003781 => D <= "11011101";	-- 0x0EC5
		when 003782 => D <= "10000010";	-- 0x0EC6
		when 003783 => D <= "10111001";	-- 0x0EC7
		when 003784 => D <= "11000010";	-- 0x0EC8
		when 003785 => D <= "10111000";	-- 0x0EC9
		when 003786 => D <= "00101110";	-- 0x0ECA
		when 003787 => D <= "11001001";	-- 0x0ECB
		when 003788 => D <= "00111110";	-- 0x0ECC
		when 003789 => D <= "00001000";	-- 0x0ECD
		when 003790 => D <= "00110010";	-- 0x0ECE
		when 003791 => D <= "11011110";	-- 0x0ECF
		when 003792 => D <= "10000010";	-- 0x0ED0
		when 003793 => D <= "00000110";	-- 0x0ED1
		when 003794 => D <= "00000001";	-- 0x0ED2
		when 003795 => D <= "11000101";	-- 0x0ED3
		when 003796 => D <= "11001101";	-- 0x0ED4
		when 003797 => D <= "10000101";	-- 0x0ED5
		when 003798 => D <= "00101110";	-- 0x0ED6
		when 003799 => D <= "00001010";	-- 0x0ED7
		when 003800 => D <= "01000111";	-- 0x0ED8
		when 003801 => D <= "00001110";	-- 0x0ED9
		when 003802 => D <= "00000000";	-- 0x0EDA
		when 003803 => D <= "00011000";	-- 0x0EDB
		when 003804 => D <= "00001111";	-- 0x0EDC
		when 003805 => D <= "00111110";	-- 0x0EDD
		when 003806 => D <= "00001000";	-- 0x0EDE
		when 003807 => D <= "00110010";	-- 0x0EDF
		when 003808 => D <= "11011110";	-- 0x0EE0
		when 003809 => D <= "10000010";	-- 0x0EE1
		when 003810 => D <= "00000110";	-- 0x0EE2
		when 003811 => D <= "00000000";	-- 0x0EE3
		when 003812 => D <= "11000101";	-- 0x0EE4
		when 003813 => D <= "11001101";	-- 0x0EE5
		when 003814 => D <= "10000101";	-- 0x0EE6
		when 003815 => D <= "00101110";	-- 0x0EE7
		when 003816 => D <= "00001010";	-- 0x0EE8
		when 003817 => D <= "01000111";	-- 0x0EE9
		when 003818 => D <= "00001110";	-- 0x0EEA
		when 003819 => D <= "00000000";	-- 0x0EEB
		when 003820 => D <= "01111000";	-- 0x0EEC
		when 003821 => D <= "10110111";	-- 0x0EED
		when 003822 => D <= "11001010";	-- 0x0EEE
		when 003823 => D <= "00000010";	-- 0x0EEF
		when 003824 => D <= "00101111";	-- 0x0EF0
		when 003825 => D <= "11011011";	-- 0x0EF1
		when 003826 => D <= "01110000";	-- 0x0EF2
		when 003827 => D <= "11100110";	-- 0x0EF3
		when 003828 => D <= "00000100";	-- 0x0EF4
		when 003829 => D <= "11001010";	-- 0x0EF5
		when 003830 => D <= "11110001";	-- 0x0EF6
		when 003831 => D <= "00101110";	-- 0x0EF7
		when 003832 => D <= "01111110";	-- 0x0EF8
		when 003833 => D <= "11010011";	-- 0x0EF9
		when 003834 => D <= "01110000";	-- 0x0EFA
		when 003835 => D <= "00100011";	-- 0x0EFB
		when 003836 => D <= "00001100";	-- 0x0EFC
		when 003837 => D <= "01111001";	-- 0x0EFD
		when 003838 => D <= "10111000";	-- 0x0EFE
		when 003839 => D <= "11000010";	-- 0x0EFF
		when 003840 => D <= "11110001";	-- 0x0F00
		when 003841 => D <= "00101110";	-- 0x0F01
		when 003842 => D <= "11001101";	-- 0x0F02
		when 003843 => D <= "11101010";	-- 0x0F03
		when 003844 => D <= "00100000";	-- 0x0F04
		when 003845 => D <= "10101111";	-- 0x0F05
		when 003846 => D <= "11010011";	-- 0x0F06
		when 003847 => D <= "01111000";	-- 0x0F07
		when 003848 => D <= "11010011";	-- 0x0F08
		when 003849 => D <= "01111001";	-- 0x0F09
		when 003850 => D <= "11011011";	-- 0x0F0A
		when 003851 => D <= "01111010";	-- 0x0F0B
		when 003852 => D <= "01100111";	-- 0x0F0C
		when 003853 => D <= "11011011";	-- 0x0F0D
		when 003854 => D <= "01111011";	-- 0x0F0E
		when 003855 => D <= "01101111";	-- 0x0F0F
		when 003856 => D <= "00010001";	-- 0x0F10
		when 003857 => D <= "00001010";	-- 0x0F11
		when 003858 => D <= "00000000";	-- 0x0F12
		when 003859 => D <= "10101111";	-- 0x0F13
		when 003860 => D <= "11101101";	-- 0x0F14
		when 003861 => D <= "01010010";	-- 0x0F15
		when 003862 => D <= "01111100";	-- 0x0F16
		when 003863 => D <= "11010011";	-- 0x0F17
		when 003864 => D <= "01111010";	-- 0x0F18
		when 003865 => D <= "01111101";	-- 0x0F19
		when 003866 => D <= "11010011";	-- 0x0F1A
		when 003867 => D <= "01111011";	-- 0x0F1B
		when 003868 => D <= "11000001";	-- 0x0F1C
		when 003869 => D <= "00000100";	-- 0x0F1D
		when 003870 => D <= "00111010";	-- 0x0F1E
		when 003871 => D <= "11011110";	-- 0x0F1F
		when 003872 => D <= "10000010";	-- 0x0F20
		when 003873 => D <= "10111000";	-- 0x0F21
		when 003874 => D <= "11000010";	-- 0x0F22
		when 003875 => D <= "11100100";	-- 0x0F23
		when 003876 => D <= "00101110";	-- 0x0F24
		when 003877 => D <= "11001001";	-- 0x0F25
		when 003878 => D <= "11111110";	-- 0x0F26
		when 003879 => D <= "00001000";	-- 0x0F27
		when 003880 => D <= "11000010";	-- 0x0F28
		when 003881 => D <= "01010011";	-- 0x0F29
		when 003882 => D <= "00101111";	-- 0x0F2A
		when 003883 => D <= "00111010";	-- 0x0F2B
		when 003884 => D <= "01001000";	-- 0x0F2C
		when 003885 => D <= "10000000";	-- 0x0F2D
		when 003886 => D <= "10110111";	-- 0x0F2E
		when 003887 => D <= "11000010";	-- 0x0F2F
		when 003888 => D <= "01001100";	-- 0x0F30
		when 003889 => D <= "00101111";	-- 0x0F31
		when 003890 => D <= "00111010";	-- 0x0F32
		when 003891 => D <= "01001001";	-- 0x0F33
		when 003892 => D <= "10000000";	-- 0x0F34
		when 003893 => D <= "10110111";	-- 0x0F35
		when 003894 => D <= "11001010";	-- 0x0F36
		when 003895 => D <= "01001001";	-- 0x0F37
		when 003896 => D <= "00101111";	-- 0x0F38
		when 003897 => D <= "00111110";	-- 0x0F39
		when 003898 => D <= "01001111";	-- 0x0F3A
		when 003899 => D <= "00110010";	-- 0x0F3B
		when 003900 => D <= "01001000";	-- 0x0F3C
		when 003901 => D <= "10000000";	-- 0x0F3D
		when 003902 => D <= "00111010";	-- 0x0F3E
		when 003903 => D <= "01001001";	-- 0x0F3F
		when 003904 => D <= "10000000";	-- 0x0F40
		when 003905 => D <= "10110111";	-- 0x0F41
		when 003906 => D <= "11001010";	-- 0x0F42
		when 003907 => D <= "01001001";	-- 0x0F43
		when 003908 => D <= "00101111";	-- 0x0F44
		when 003909 => D <= "00111101";	-- 0x0F45
		when 003910 => D <= "00110010";	-- 0x0F46
		when 003911 => D <= "01001001";	-- 0x0F47
		when 003912 => D <= "10000000";	-- 0x0F48
		when 003913 => D <= "11000011";	-- 0x0F49
		when 003914 => D <= "01010000";	-- 0x0F4A
		when 003915 => D <= "00101111";	-- 0x0F4B
		when 003916 => D <= "00111101";	-- 0x0F4C
		when 003917 => D <= "00110010";	-- 0x0F4D
		when 003918 => D <= "01001000";	-- 0x0F4E
		when 003919 => D <= "10000000";	-- 0x0F4F
		when 003920 => D <= "11000011";	-- 0x0F50
		when 003921 => D <= "11111100";	-- 0x0F51
		when 003922 => D <= "00101111";	-- 0x0F52
		when 003923 => D <= "11111110";	-- 0x0F53
		when 003924 => D <= "00011010";	-- 0x0F54
		when 003925 => D <= "11000010";	-- 0x0F55
		when 003926 => D <= "01011110";	-- 0x0F56
		when 003927 => D <= "00101111";	-- 0x0F57
		when 003928 => D <= "11001101";	-- 0x0F58
		when 003929 => D <= "00010001";	-- 0x0F59
		when 003930 => D <= "00100001";	-- 0x0F5A
		when 003931 => D <= "11000011";	-- 0x0F5B
		when 003932 => D <= "11111100";	-- 0x0F5C
		when 003933 => D <= "00101111";	-- 0x0F5D
		when 003934 => D <= "11111110";	-- 0x0F5E
		when 003935 => D <= "00011110";	-- 0x0F5F
		when 003936 => D <= "11000010";	-- 0x0F60
		when 003937 => D <= "01101101";	-- 0x0F61
		when 003938 => D <= "00101111";	-- 0x0F62
		when 003939 => D <= "10101111";	-- 0x0F63
		when 003940 => D <= "00110010";	-- 0x0F64
		when 003941 => D <= "01001000";	-- 0x0F65
		when 003942 => D <= "10000000";	-- 0x0F66
		when 003943 => D <= "00110010";	-- 0x0F67
		when 003944 => D <= "01001001";	-- 0x0F68
		when 003945 => D <= "10000000";	-- 0x0F69
		when 003946 => D <= "11000011";	-- 0x0F6A
		when 003947 => D <= "11111100";	-- 0x0F6B
		when 003948 => D <= "00101111";	-- 0x0F6C
		when 003949 => D <= "11111110";	-- 0x0F6D
		when 003950 => D <= "00001011";	-- 0x0F6E
		when 003951 => D <= "11000010";	-- 0x0F6F
		when 003952 => D <= "10000000";	-- 0x0F70
		when 003953 => D <= "00101111";	-- 0x0F71
		when 003954 => D <= "00111010";	-- 0x0F72
		when 003955 => D <= "01001001";	-- 0x0F73
		when 003956 => D <= "10000000";	-- 0x0F74
		when 003957 => D <= "10110111";	-- 0x0F75
		when 003958 => D <= "11001010";	-- 0x0F76
		when 003959 => D <= "01111101";	-- 0x0F77
		when 003960 => D <= "00101111";	-- 0x0F78
		when 003961 => D <= "00111101";	-- 0x0F79
		when 003962 => D <= "00110010";	-- 0x0F7A
		when 003963 => D <= "01001001";	-- 0x0F7B
		when 003964 => D <= "10000000";	-- 0x0F7C
		when 003965 => D <= "11000011";	-- 0x0F7D
		when 003966 => D <= "11111100";	-- 0x0F7E
		when 003967 => D <= "00101111";	-- 0x0F7F
		when 003968 => D <= "11111110";	-- 0x0F80
		when 003969 => D <= "00001010";	-- 0x0F81
		when 003970 => D <= "11000010";	-- 0x0F82
		when 003971 => D <= "10011010";	-- 0x0F83
		when 003972 => D <= "00101111";	-- 0x0F84
		when 003973 => D <= "00111010";	-- 0x0F85
		when 003974 => D <= "01001001";	-- 0x0F86
		when 003975 => D <= "10000000";	-- 0x0F87
		when 003976 => D <= "11111110";	-- 0x0F88
		when 003977 => D <= "00000111";	-- 0x0F89
		when 003978 => D <= "11010010";	-- 0x0F8A
		when 003979 => D <= "10010100";	-- 0x0F8B
		when 003980 => D <= "00101111";	-- 0x0F8C
		when 003981 => D <= "00111100";	-- 0x0F8D
		when 003982 => D <= "00110010";	-- 0x0F8E
		when 003983 => D <= "01001001";	-- 0x0F8F
		when 003984 => D <= "10000000";	-- 0x0F90
		when 003985 => D <= "11000011";	-- 0x0F91
		when 003986 => D <= "10010111";	-- 0x0F92
		when 003987 => D <= "00101111";	-- 0x0F93
		when 003988 => D <= "11001101";	-- 0x0F94
		when 003989 => D <= "00110000";	-- 0x0F95
		when 003990 => D <= "00101101";	-- 0x0F96
		when 003991 => D <= "11000011";	-- 0x0F97
		when 003992 => D <= "11111100";	-- 0x0F98
		when 003993 => D <= "00101111";	-- 0x0F99
		when 003994 => D <= "11111110";	-- 0x0F9A
		when 003995 => D <= "00001001";	-- 0x0F9B
		when 003996 => D <= "11000010";	-- 0x0F9C
		when 003997 => D <= "11000111";	-- 0x0F9D
		when 003998 => D <= "00101111";	-- 0x0F9E
		when 003999 => D <= "00111010";	-- 0x0F9F
		when 004000 => D <= "01001000";	-- 0x0FA0
		when 004001 => D <= "10000000";	-- 0x0FA1
		when 004002 => D <= "11111110";	-- 0x0FA2
		when 004003 => D <= "01001111";	-- 0x0FA3
		when 004004 => D <= "11000010";	-- 0x0FA4
		when 004005 => D <= "11000000";	-- 0x0FA5
		when 004006 => D <= "00101111";	-- 0x0FA6
		when 004007 => D <= "10101111";	-- 0x0FA7
		when 004008 => D <= "00110010";	-- 0x0FA8
		when 004009 => D <= "01001000";	-- 0x0FA9
		when 004010 => D <= "10000000";	-- 0x0FAA
		when 004011 => D <= "00111010";	-- 0x0FAB
		when 004012 => D <= "01001001";	-- 0x0FAC
		when 004013 => D <= "10000000";	-- 0x0FAD
		when 004014 => D <= "11111110";	-- 0x0FAE
		when 004015 => D <= "00000111";	-- 0x0FAF
		when 004016 => D <= "11000010";	-- 0x0FB0
		when 004017 => D <= "10111001";	-- 0x0FB1
		when 004018 => D <= "00101111";	-- 0x0FB2
		when 004019 => D <= "11001101";	-- 0x0FB3
		when 004020 => D <= "00110000";	-- 0x0FB4
		when 004021 => D <= "00101101";	-- 0x0FB5
		when 004022 => D <= "11000011";	-- 0x0FB6
		when 004023 => D <= "10111101";	-- 0x0FB7
		when 004024 => D <= "00101111";	-- 0x0FB8
		when 004025 => D <= "00111100";	-- 0x0FB9
		when 004026 => D <= "00110010";	-- 0x0FBA
		when 004027 => D <= "01001001";	-- 0x0FBB
		when 004028 => D <= "10000000";	-- 0x0FBC
		when 004029 => D <= "11000011";	-- 0x0FBD
		when 004030 => D <= "11000100";	-- 0x0FBE
		when 004031 => D <= "00101111";	-- 0x0FBF
		when 004032 => D <= "00111100";	-- 0x0FC0
		when 004033 => D <= "00110010";	-- 0x0FC1
		when 004034 => D <= "01001000";	-- 0x0FC2
		when 004035 => D <= "10000000";	-- 0x0FC3
		when 004036 => D <= "11000011";	-- 0x0FC4
		when 004037 => D <= "11111100";	-- 0x0FC5
		when 004038 => D <= "00101111";	-- 0x0FC6
		when 004039 => D <= "11111110";	-- 0x0FC7
		when 004040 => D <= "00001101";	-- 0x0FC8
		when 004041 => D <= "11000010";	-- 0x0FC9
		when 004042 => D <= "11010011";	-- 0x0FCA
		when 004043 => D <= "00101111";	-- 0x0FCB
		when 004044 => D <= "10101111";	-- 0x0FCC
		when 004045 => D <= "00110010";	-- 0x0FCD
		when 004046 => D <= "01001000";	-- 0x0FCE
		when 004047 => D <= "10000000";	-- 0x0FCF
		when 004048 => D <= "11000011";	-- 0x0FD0
		when 004049 => D <= "11111100";	-- 0x0FD1
		when 004050 => D <= "00101111";	-- 0x0FD2
		when 004051 => D <= "11111110";	-- 0x0FD3
		when 004052 => D <= "00010110";	-- 0x0FD4
		when 004053 => D <= "11000010";	-- 0x0FD5
		when 004054 => D <= "11011110";	-- 0x0FD6
		when 004055 => D <= "00101111";	-- 0x0FD7
		when 004056 => D <= "11001101";	-- 0x0FD8
		when 004057 => D <= "10101011";	-- 0x0FD9
		when 004058 => D <= "00101101";	-- 0x0FDA
		when 004059 => D <= "11000011";	-- 0x0FDB
		when 004060 => D <= "11111100";	-- 0x0FDC
		when 004061 => D <= "00101111";	-- 0x0FDD
		when 004062 => D <= "11111110";	-- 0x0FDE
		when 004063 => D <= "01111111";	-- 0x0FDF
		when 004064 => D <= "11000010";	-- 0x0FE0
		when 004065 => D <= "11110100";	-- 0x0FE1
		when 004066 => D <= "00101111";	-- 0x0FE2
		when 004067 => D <= "00111010";	-- 0x0FE3
		when 004068 => D <= "01001000";	-- 0x0FE4
		when 004069 => D <= "10000000";	-- 0x0FE5
		when 004070 => D <= "10110111";	-- 0x0FE6
		when 004071 => D <= "11001010";	-- 0x0FE7
		when 004072 => D <= "11110001";	-- 0x0FE8
		when 004073 => D <= "00101111";	-- 0x0FE9
		when 004074 => D <= "00111101";	-- 0x0FEA
		when 004075 => D <= "00110010";	-- 0x0FEB
		when 004076 => D <= "01001000";	-- 0x0FEC
		when 004077 => D <= "10000000";	-- 0x0FED
		when 004078 => D <= "11001101";	-- 0x0FEE
		when 004079 => D <= "00010010";	-- 0x0FEF
		when 004080 => D <= "00101110";	-- 0x0FF0
		when 004081 => D <= "11000011";	-- 0x0FF1
		when 004082 => D <= "11111100";	-- 0x0FF2
		when 004083 => D <= "00101111";	-- 0x0FF3
		when 004084 => D <= "11111110";	-- 0x0FF4
		when 004085 => D <= "00000111";	-- 0x0FF5
		when 004086 => D <= "11000010";	-- 0x0FF6
		when 004087 => D <= "11111100";	-- 0x0FF7
		when 004088 => D <= "00101111";	-- 0x0FF8
		when 004089 => D <= "11001101";	-- 0x0FF9
		when 004090 => D <= "00010010";	-- 0x0FFA
		when 004091 => D <= "00101110";	-- 0x0FFB
		when 004092 => D <= "11001001";	-- 0x0FFC
		when 004093 => D <= "11100110";	-- 0x0FFD
		when 004094 => D <= "01111111";	-- 0x0FFE
		when 004095 => D <= "11110101";	-- 0x0FFF
		when 004096 => D <= "10101111";	-- 0x1000
		when 004097 => D <= "00110010";	-- 0x1001
		when 004098 => D <= "01000110";	-- 0x1002
		when 004099 => D <= "10000000";	-- 0x1003
		when 004100 => D <= "11001101";	-- 0x1004
		when 004101 => D <= "01011000";	-- 0x1005
		when 004102 => D <= "00100001";	-- 0x1006
		when 004103 => D <= "11001101";	-- 0x1007
		when 004104 => D <= "10010100";	-- 0x1008
		when 004105 => D <= "00101100";	-- 0x1009
		when 004106 => D <= "11001101";	-- 0x100A
		when 004107 => D <= "10111101";	-- 0x100B
		when 004108 => D <= "00101100";	-- 0x100C
		when 004109 => D <= "00001010";	-- 0x100D
		when 004110 => D <= "01011111";	-- 0x100E
		when 004111 => D <= "00111010";	-- 0x100F
		when 004112 => D <= "01001000";	-- 0x1010
		when 004113 => D <= "10000000";	-- 0x1011
		when 004114 => D <= "00111100";	-- 0x1012
		when 004115 => D <= "10111011";	-- 0x1013
		when 004116 => D <= "11001010";	-- 0x1014
		when 004117 => D <= "00011011";	-- 0x1015
		when 004118 => D <= "00110000";	-- 0x1016
		when 004119 => D <= "11011010";	-- 0x1017
		when 004120 => D <= "00011011";	-- 0x1018
		when 004121 => D <= "00110000";	-- 0x1019
		when 004122 => D <= "00000010";	-- 0x101A
		when 004123 => D <= "01111110";	-- 0x101B
		when 004124 => D <= "00110010";	-- 0x101C
		when 004125 => D <= "11011100";	-- 0x101D
		when 004126 => D <= "10000010";	-- 0x101E
		when 004127 => D <= "11111110";	-- 0x101F
		when 004128 => D <= "00100000";	-- 0x1020
		when 004129 => D <= "11001010";	-- 0x1021
		when 004130 => D <= "00101111";	-- 0x1022
		when 004131 => D <= "00110000";	-- 0x1023
		when 004132 => D <= "11001101";	-- 0x1024
		when 004133 => D <= "01000110";	-- 0x1025
		when 004134 => D <= "00100010";	-- 0x1026
		when 004135 => D <= "00111110";	-- 0x1027
		when 004136 => D <= "00001010";	-- 0x1028
		when 004137 => D <= "11001101";	-- 0x1029
		when 004138 => D <= "11110011";	-- 0x102A
		when 004139 => D <= "00100000";	-- 0x102B
		when 004140 => D <= "11001101";	-- 0x102C
		when 004141 => D <= "10010100";	-- 0x102D
		when 004142 => D <= "00101100";	-- 0x102E
		when 004143 => D <= "11001101";	-- 0x102F
		when 004144 => D <= "01000010";	-- 0x1030
		when 004145 => D <= "00100010";	-- 0x1031
		when 004146 => D <= "11110001";	-- 0x1032
		when 004147 => D <= "11110101";	-- 0x1033
		when 004148 => D <= "01110111";	-- 0x1034
		when 004149 => D <= "10110111";	-- 0x1035
		when 004150 => D <= "11001101";	-- 0x1036
		when 004151 => D <= "11110011";	-- 0x1037
		when 004152 => D <= "00100000";	-- 0x1038
		when 004153 => D <= "00111110";	-- 0x1039
		when 004154 => D <= "00000001";	-- 0x103A
		when 004155 => D <= "00110010";	-- 0x103B
		when 004156 => D <= "01000110";	-- 0x103C
		when 004157 => D <= "10000000";	-- 0x103D
		when 004158 => D <= "11001101";	-- 0x103E
		when 004159 => D <= "01011000";	-- 0x103F
		when 004160 => D <= "00100001";	-- 0x1040
		when 004161 => D <= "11001101";	-- 0x1041
		when 004162 => D <= "10010100";	-- 0x1042
		when 004163 => D <= "00101100";	-- 0x1043
		when 004164 => D <= "00111010";	-- 0x1044
		when 004165 => D <= "11011100";	-- 0x1045
		when 004166 => D <= "10000010";	-- 0x1046
		when 004167 => D <= "11111110";	-- 0x1047
		when 004168 => D <= "00100000";	-- 0x1048
		when 004169 => D <= "11001010";	-- 0x1049
		when 004170 => D <= "01011010";	-- 0x104A
		when 004171 => D <= "00110000";	-- 0x104B
		when 004172 => D <= "11001101";	-- 0x104C
		when 004173 => D <= "01000110";	-- 0x104D
		when 004174 => D <= "00100010";	-- 0x104E
		when 004175 => D <= "00111110";	-- 0x104F
		when 004176 => D <= "00001010";	-- 0x1050
		when 004177 => D <= "11001101";	-- 0x1051
		when 004178 => D <= "11110011";	-- 0x1052
		when 004179 => D <= "00100000";	-- 0x1053
		when 004180 => D <= "11001101";	-- 0x1054
		when 004181 => D <= "10010100";	-- 0x1055
		when 004182 => D <= "00101100";	-- 0x1056
		when 004183 => D <= "11001101";	-- 0x1057
		when 004184 => D <= "01000010";	-- 0x1058
		when 004185 => D <= "00100010";	-- 0x1059
		when 004186 => D <= "11110001";	-- 0x105A
		when 004187 => D <= "11001101";	-- 0x105B
		when 004188 => D <= "11110011";	-- 0x105C
		when 004189 => D <= "00100000";	-- 0x105D
		when 004190 => D <= "00111010";	-- 0x105E
		when 004191 => D <= "01001000";	-- 0x105F
		when 004192 => D <= "10000000";	-- 0x1060
		when 004193 => D <= "00111100";	-- 0x1061
		when 004194 => D <= "00110010";	-- 0x1062
		when 004195 => D <= "01001000";	-- 0x1063
		when 004196 => D <= "10000000";	-- 0x1064
		when 004197 => D <= "11111110";	-- 0x1065
		when 004198 => D <= "01001111";	-- 0x1066
		when 004199 => D <= "11001010";	-- 0x1067
		when 004200 => D <= "10001000";	-- 0x1068
		when 004201 => D <= "00110000";	-- 0x1069
		when 004202 => D <= "11011010";	-- 0x106A
		when 004203 => D <= "10001000";	-- 0x106B
		when 004204 => D <= "00110000";	-- 0x106C
		when 004205 => D <= "10101111";	-- 0x106D
		when 004206 => D <= "00110010";	-- 0x106E
		when 004207 => D <= "01001000";	-- 0x106F
		when 004208 => D <= "10000000";	-- 0x1070
		when 004209 => D <= "00111010";	-- 0x1071
		when 004210 => D <= "01001001";	-- 0x1072
		when 004211 => D <= "10000000";	-- 0x1073
		when 004212 => D <= "00111100";	-- 0x1074
		when 004213 => D <= "00110010";	-- 0x1075
		when 004214 => D <= "01001001";	-- 0x1076
		when 004215 => D <= "10000000";	-- 0x1077
		when 004216 => D <= "11111110";	-- 0x1078
		when 004217 => D <= "00000111";	-- 0x1079
		when 004218 => D <= "11001010";	-- 0x107A
		when 004219 => D <= "10001000";	-- 0x107B
		when 004220 => D <= "00110000";	-- 0x107C
		when 004221 => D <= "11011010";	-- 0x107D
		when 004222 => D <= "10001000";	-- 0x107E
		when 004223 => D <= "00110000";	-- 0x107F
		when 004224 => D <= "00111110";	-- 0x1080
		when 004225 => D <= "00000111";	-- 0x1081
		when 004226 => D <= "00110010";	-- 0x1082
		when 004227 => D <= "01001001";	-- 0x1083
		when 004228 => D <= "10000000";	-- 0x1084
		when 004229 => D <= "11001101";	-- 0x1085
		when 004230 => D <= "00110000";	-- 0x1086
		when 004231 => D <= "00101101";	-- 0x1087
		when 004232 => D <= "11001001";	-- 0x1088
		when 004233 => D <= "11001101";	-- 0x1089
		when 004234 => D <= "00001000";	-- 0x108A
		when 004235 => D <= "00100000";	-- 0x108B
		when 004236 => D <= "11001010";	-- 0x108C
		when 004237 => D <= "10110110";	-- 0x108D
		when 004238 => D <= "00110000";	-- 0x108E
		when 004239 => D <= "10101111";	-- 0x108F
		when 004240 => D <= "00110010";	-- 0x1090
		when 004241 => D <= "00010110";	-- 0x1091
		when 004242 => D <= "10000000";	-- 0x1092
		when 004243 => D <= "11001101";	-- 0x1093
		when 004244 => D <= "00101001";	-- 0x1094
		when 004245 => D <= "00100000";	-- 0x1095
		when 004246 => D <= "11111110";	-- 0x1096
		when 004247 => D <= "00010011";	-- 0x1097
		when 004248 => D <= "11000010";	-- 0x1098
		when 004249 => D <= "10101110";	-- 0x1099
		when 004250 => D <= "00110000";	-- 0x109A
		when 004251 => D <= "11001101";	-- 0x109B
		when 004252 => D <= "00101001";	-- 0x109C
		when 004253 => D <= "00100000";	-- 0x109D
		when 004254 => D <= "11111110";	-- 0x109E
		when 004255 => D <= "00000011";	-- 0x109F
		when 004256 => D <= "11000010";	-- 0x10A0
		when 004257 => D <= "10100110";	-- 0x10A1
		when 004258 => D <= "00110000";	-- 0x10A2
		when 004259 => D <= "11000011";	-- 0x10A3
		when 004260 => D <= "10011010";	-- 0x10A4
		when 004261 => D <= "00111111";	-- 0x10A5
		when 004262 => D <= "11111110";	-- 0x10A6
		when 004263 => D <= "00010001";	-- 0x10A7
		when 004264 => D <= "11000010";	-- 0x10A8
		when 004265 => D <= "10011011";	-- 0x10A9
		when 004266 => D <= "00110000";	-- 0x10AA
		when 004267 => D <= "11000011";	-- 0x10AB
		when 004268 => D <= "10110110";	-- 0x10AC
		when 004269 => D <= "00110000";	-- 0x10AD
		when 004270 => D <= "00110010";	-- 0x10AE
		when 004271 => D <= "00010111";	-- 0x10AF
		when 004272 => D <= "10000000";	-- 0x10B0
		when 004273 => D <= "00111110";	-- 0x10B1
		when 004274 => D <= "11111111";	-- 0x10B2
		when 004275 => D <= "00110010";	-- 0x10B3
		when 004276 => D <= "00010110";	-- 0x10B4
		when 004277 => D <= "10000000";	-- 0x10B5
		when 004278 => D <= "11001001";	-- 0x10B6
		when 004279 => D <= "11001101";	-- 0x10B7
		when 004280 => D <= "10001001";	-- 0x10B8
		when 004281 => D <= "00110000";	-- 0x10B9
		when 004282 => D <= "11111101";	-- 0x10BA
		when 004283 => D <= "11100101";	-- 0x10BB
		when 004284 => D <= "11011101";	-- 0x10BC
		when 004285 => D <= "11100101";	-- 0x10BD
		when 004286 => D <= "11100101";	-- 0x10BE
		when 004287 => D <= "11010101";	-- 0x10BF
		when 004288 => D <= "11000101";	-- 0x10C0
		when 004289 => D <= "00111010";	-- 0x10C1
		when 004290 => D <= "00000100";	-- 0x10C2
		when 004291 => D <= "10000000";	-- 0x10C3
		when 004292 => D <= "11111110";	-- 0x10C4
		when 004293 => D <= "00000001";	-- 0x10C5
		when 004294 => D <= "11000010";	-- 0x10C6
		when 004295 => D <= "11010000";	-- 0x10C7
		when 004296 => D <= "00110000";	-- 0x10C8
		when 004297 => D <= "11000101";	-- 0x10C9
		when 004298 => D <= "11001011";	-- 0x10CA
		when 004299 => D <= "10111001";	-- 0x10CB
		when 004300 => D <= "11001101";	-- 0x10CC
		when 004301 => D <= "11011001";	-- 0x10CD
		when 004302 => D <= "00100000";	-- 0x10CE
		when 004303 => D <= "11000001";	-- 0x10CF
		when 004304 => D <= "01111001";	-- 0x10D0
		when 004305 => D <= "11100110";	-- 0x10D1
		when 004306 => D <= "01111111";	-- 0x10D2
		when 004307 => D <= "11111110";	-- 0x10D3
		when 004308 => D <= "00100000";	-- 0x10D4
		when 004309 => D <= "11011010";	-- 0x10D5
		when 004310 => D <= "11011101";	-- 0x10D6
		when 004311 => D <= "00110000";	-- 0x10D7
		when 004312 => D <= "11111110";	-- 0x10D8
		when 004313 => D <= "01111111";	-- 0x10D9
		when 004314 => D <= "11000010";	-- 0x10DA
		when 004315 => D <= "11100011";	-- 0x10DB
		when 004316 => D <= "00110000";	-- 0x10DC
		when 004317 => D <= "11001101";	-- 0x10DD
		when 004318 => D <= "00100110";	-- 0x10DE
		when 004319 => D <= "00101111";	-- 0x10DF
		when 004320 => D <= "11000011";	-- 0x10E0
		when 004321 => D <= "11100110";	-- 0x10E1
		when 004322 => D <= "00110000";	-- 0x10E2
		when 004323 => D <= "11001101";	-- 0x10E3
		when 004324 => D <= "11111101";	-- 0x10E4
		when 004325 => D <= "00101111";	-- 0x10E5
		when 004326 => D <= "11000001";	-- 0x10E6
		when 004327 => D <= "11010001";	-- 0x10E7
		when 004328 => D <= "11100001";	-- 0x10E8
		when 004329 => D <= "11011101";	-- 0x10E9
		when 004330 => D <= "11100001";	-- 0x10EA
		when 004331 => D <= "11111101";	-- 0x10EB
		when 004332 => D <= "11100001";	-- 0x10EC
		when 004333 => D <= "01111001";	-- 0x10ED
		when 004334 => D <= "11001001";	-- 0x10EE
		when 004335 => D <= "00001110";	-- 0x10EF
		when 004336 => D <= "00001101";	-- 0x10F0
		when 004337 => D <= "11001101";	-- 0x10F1
		when 004338 => D <= "10110111";	-- 0x10F2
		when 004339 => D <= "00110000";	-- 0x10F3
		when 004340 => D <= "00001110";	-- 0x10F4
		when 004341 => D <= "00001010";	-- 0x10F5
		when 004342 => D <= "11000011";	-- 0x10F6
		when 004343 => D <= "10110111";	-- 0x10F7
		when 004344 => D <= "00110000";	-- 0x10F8
		when 004345 => D <= "11001101";	-- 0x10F9
		when 004346 => D <= "00101001";	-- 0x10FA
		when 004347 => D <= "00100000";	-- 0x10FB
		when 004348 => D <= "01001111";	-- 0x10FC
		when 004349 => D <= "11001101";	-- 0x10FD
		when 004350 => D <= "10110111";	-- 0x10FE
		when 004351 => D <= "00110000";	-- 0x10FF
		when 004352 => D <= "11111110";	-- 0x1100
		when 004353 => D <= "00001101";	-- 0x1101
		when 004354 => D <= "11000010";	-- 0x1102
		when 004355 => D <= "11111001";	-- 0x1103
		when 004356 => D <= "00110000";	-- 0x1104
		when 004357 => D <= "00111010";	-- 0x1105
		when 004358 => D <= "01001001";	-- 0x1106
		when 004359 => D <= "10000000";	-- 0x1107
		when 004360 => D <= "01000111";	-- 0x1108
		when 004361 => D <= "11001101";	-- 0x1109
		when 004362 => D <= "10000101";	-- 0x110A
		when 004363 => D <= "00101110";	-- 0x110B
		when 004364 => D <= "11011101";	-- 0x110C
		when 004365 => D <= "00100001";	-- 0x110D
		when 004366 => D <= "11101111";	-- 0x110E
		when 004367 => D <= "10000010";	-- 0x110F
		when 004368 => D <= "00001010";	-- 0x1110
		when 004369 => D <= "10110111";	-- 0x1111
		when 004370 => D <= "11001010";	-- 0x1112
		when 004371 => D <= "00100000";	-- 0x1113
		when 004372 => D <= "00110001";	-- 0x1114
		when 004373 => D <= "01000110";	-- 0x1115
		when 004374 => D <= "11011101";	-- 0x1116
		when 004375 => D <= "01110000";	-- 0x1117
		when 004376 => D <= "00000000";	-- 0x1118
		when 004377 => D <= "00100011";	-- 0x1119
		when 004378 => D <= "11011101";	-- 0x111A
		when 004379 => D <= "00100011";	-- 0x111B
		when 004380 => D <= "00111101";	-- 0x111C
		when 004381 => D <= "11000011";	-- 0x111D
		when 004382 => D <= "00010001";	-- 0x111E
		when 004383 => D <= "00110001";	-- 0x111F
		when 004384 => D <= "11011101";	-- 0x1120
		when 004385 => D <= "00110110";	-- 0x1121
		when 004386 => D <= "00000000";	-- 0x1122
		when 004387 => D <= "00000000";	-- 0x1123
		when 004388 => D <= "00100001";	-- 0x1124
		when 004389 => D <= "11101111";	-- 0x1125
		when 004390 => D <= "10000010";	-- 0x1126
		when 004391 => D <= "11001101";	-- 0x1127
		when 004392 => D <= "11101111";	-- 0x1128
		when 004393 => D <= "00110000";	-- 0x1129
		when 004394 => D <= "11001001";	-- 0x112A
		when 004395 => D <= "10000101";	-- 0x112B
		when 004396 => D <= "00110011";	-- 0x112C
		when 004397 => D <= "10010010";	-- 0x112D
		when 004398 => D <= "00110011";	-- 0x112E
		when 004399 => D <= "10100110";	-- 0x112F
		when 004400 => D <= "00110011";	-- 0x1130
		when 004401 => D <= "10110000";	-- 0x1131
		when 004402 => D <= "00110011";	-- 0x1132
		when 004403 => D <= "11111101";	-- 0x1133
		when 004404 => D <= "00110011";	-- 0x1134
		when 004405 => D <= "00000001";	-- 0x1135
		when 004406 => D <= "00110100";	-- 0x1136
		when 004407 => D <= "00000101";	-- 0x1137
		when 004408 => D <= "00110100";	-- 0x1138
		when 004409 => D <= "00001001";	-- 0x1139
		when 004410 => D <= "00110100";	-- 0x113A
		when 004411 => D <= "11001000";	-- 0x113B
		when 004412 => D <= "00110100";	-- 0x113C
		when 004413 => D <= "11100101";	-- 0x113D
		when 004414 => D <= "00110101";	-- 0x113E
		when 004415 => D <= "11111000";	-- 0x113F
		when 004416 => D <= "00110101";	-- 0x1140
		when 004417 => D <= "01110111";	-- 0x1141
		when 004418 => D <= "00110111";	-- 0x1142
		when 004419 => D <= "11011100";	-- 0x1143
		when 004420 => D <= "00110111";	-- 0x1144
		when 004421 => D <= "01011101";	-- 0x1145
		when 004422 => D <= "00111000";	-- 0x1146
		when 004423 => D <= "10000010";	-- 0x1147
		when 004424 => D <= "00111000";	-- 0x1148
		when 004425 => D <= "10111111";	-- 0x1149
		when 004426 => D <= "00111000";	-- 0x114A
		when 004427 => D <= "11100001";	-- 0x114B
		when 004428 => D <= "00111000";	-- 0x114C
		when 004429 => D <= "11101010";	-- 0x114D
		when 004430 => D <= "00111000";	-- 0x114E
		when 004431 => D <= "00001100";	-- 0x114F
		when 004432 => D <= "00111010";	-- 0x1150
		when 004433 => D <= "01001110";	-- 0x1151
		when 004434 => D <= "00111001";	-- 0x1152
		when 004435 => D <= "11100110";	-- 0x1153
		when 004436 => D <= "00111010";	-- 0x1154
		when 004437 => D <= "10011001";	-- 0x1155
		when 004438 => D <= "00111011";	-- 0x1156
		when 004439 => D <= "00001011";	-- 0x1157
		when 004440 => D <= "00111100";	-- 0x1158
		when 004441 => D <= "10011100";	-- 0x1159
		when 004442 => D <= "00110011";	-- 0x115A
		when 004443 => D <= "11101111";	-- 0x115B
		when 004444 => D <= "00110111";	-- 0x115C
		when 004445 => D <= "01100100";	-- 0x115D
		when 004446 => D <= "00111000";	-- 0x115E
		when 004447 => D <= "01101111";	-- 0x115F
		when 004448 => D <= "00111000";	-- 0x1160
		when 004449 => D <= "10111101";	-- 0x1161
		when 004450 => D <= "00110011";	-- 0x1162
		when 004451 => D <= "11100010";	-- 0x1163
		when 004452 => D <= "00110011";	-- 0x1164
		when 004453 => D <= "01111111";	-- 0x1165
		when 004454 => D <= "00110110";	-- 0x1166
		when 004455 => D <= "10010100";	-- 0x1167
		when 004456 => D <= "00110110";	-- 0x1168
		when 004457 => D <= "10101011";	-- 0x1169
		when 004458 => D <= "00110110";	-- 0x116A
		when 004459 => D <= "00010110";	-- 0x116B
		when 004460 => D <= "00110111";	-- 0x116C
		when 004461 => D <= "00001101";	-- 0x116D
		when 004462 => D <= "00110111";	-- 0x116E
		when 004463 => D <= "00010011";	-- 0x116F
		when 004464 => D <= "00110111";	-- 0x1170
		when 004465 => D <= "11000010";	-- 0x1171
		when 004466 => D <= "00110110";	-- 0x1172
		when 004467 => D <= "00011011";	-- 0x1173
		when 004468 => D <= "00111001";	-- 0x1174
		when 004469 => D <= "00010010";	-- 0x1175
		when 004470 => D <= "00111001";	-- 0x1176
		when 004471 => D <= "10011011";	-- 0x1177
		when 004472 => D <= "00111000";	-- 0x1178
		when 004473 => D <= "10101101";	-- 0x1179
		when 004474 => D <= "00111000";	-- 0x117A
		when 004475 => D <= "00100010";	-- 0x117B
		when 004476 => D <= "00111001";	-- 0x117C
		when 004477 => D <= "00111101";	-- 0x117D
		when 004478 => D <= "00111001";	-- 0x117E
		when 004479 => D <= "11101110";	-- 0x117F
		when 004480 => D <= "00111000";	-- 0x1180
		when 004481 => D <= "00001000";	-- 0x1181
		when 004482 => D <= "00111010";	-- 0x1182
		when 004483 => D <= "11111100";	-- 0x1183
		when 004484 => D <= "00111011";	-- 0x1184
		when 004485 => D <= "00001000";	-- 0x1185
		when 004486 => D <= "00111100";	-- 0x1186
		when 004487 => D <= "01010110";	-- 0x1187
		when 004488 => D <= "11010111";	-- 0x1188
		when 004489 => D <= "10000010";	-- 0x1189
		when 004490 => D <= "00000000";	-- 0x118A
		when 004491 => D <= "00000010";	-- 0x118B
		when 004492 => D <= "01010010";	-- 0x118C
		when 004493 => D <= "11010111";	-- 0x118D
		when 004494 => D <= "10000001";	-- 0x118E
		when 004495 => D <= "00000000";	-- 0x118F
		when 004496 => D <= "00000010";	-- 0x1190
		when 004497 => D <= "01001100";	-- 0x1191
		when 004498 => D <= "11001001";	-- 0x1192
		when 004499 => D <= "10000011";	-- 0x1193
		when 004500 => D <= "00000000";	-- 0x1194
		when 004501 => D <= "00000010";	-- 0x1195
		when 004502 => D <= "01010010";	-- 0x1196
		when 004503 => D <= "11000101";	-- 0x1197
		when 004504 => D <= "10000100";	-- 0x1198
		when 004505 => D <= "00000000";	-- 0x1199
		when 004506 => D <= "00000010";	-- 0x119A
		when 004507 => D <= "01010111";	-- 0x119B
		when 004508 => D <= "01000101";	-- 0x119C
		when 004509 => D <= "01001110";	-- 0x119D
		when 004510 => D <= "11001110";	-- 0x119E
		when 004511 => D <= "10001011";	-- 0x119F
		when 004512 => D <= "00000000";	-- 0x11A0
		when 004513 => D <= "00000010";	-- 0x11A1
		when 004514 => D <= "01010111";	-- 0x11A2
		when 004515 => D <= "11001000";	-- 0x11A3
		when 004516 => D <= "10001100";	-- 0x11A4
		when 004517 => D <= "00000000";	-- 0x11A5
		when 004518 => D <= "00000010";	-- 0x11A6
		when 004519 => D <= "01010010";	-- 0x11A7
		when 004520 => D <= "11001011";	-- 0x11A8
		when 004521 => D <= "10001101";	-- 0x11A9
		when 004522 => D <= "00000000";	-- 0x11AA
		when 004523 => D <= "00000010";	-- 0x11AB
		when 004524 => D <= "01010011";	-- 0x11AC
		when 004525 => D <= "01000101";	-- 0x11AD
		when 004526 => D <= "01010100";	-- 0x11AE
		when 004527 => D <= "01011010";	-- 0x11AF
		when 004528 => D <= "11000101";	-- 0x11B0
		when 004529 => D <= "10010110";	-- 0x11B1
		when 004530 => D <= "00000000";	-- 0x11B2
		when 004531 => D <= "00000010";	-- 0x11B3
		when 004532 => D <= "01000101";	-- 0x11B4
		when 004533 => D <= "01001110";	-- 0x11B5
		when 004534 => D <= "01000100";	-- 0x11B6
		when 004535 => D <= "11000101";	-- 0x11B7
		when 004536 => D <= "10001010";	-- 0x11B8
		when 004537 => D <= "00000000";	-- 0x11B9
		when 004538 => D <= "00000010";	-- 0x11BA
		when 004539 => D <= "01010000";	-- 0x11BB
		when 004540 => D <= "01001111";	-- 0x11BC
		when 004541 => D <= "01010010";	-- 0x11BD
		when 004542 => D <= "11010100";	-- 0x11BE
		when 004543 => D <= "10011011";	-- 0x11BF
		when 004544 => D <= "00000000";	-- 0x11C0
		when 004545 => D <= "00000010";	-- 0x11C1
		when 004546 => D <= "01010011";	-- 0x11C2
		when 004547 => D <= "11001111";	-- 0x11C3
		when 004548 => D <= "10100100";	-- 0x11C4
		when 004549 => D <= "00000000";	-- 0x11C5
		when 004550 => D <= "00000010";	-- 0x11C6
		when 004551 => D <= "01010111";	-- 0x11C7
		when 004552 => D <= "01001001";	-- 0x11C8
		when 004553 => D <= "01000101";	-- 0x11C9
		when 004554 => D <= "01000100";	-- 0x11CA
		when 004555 => D <= "01000101";	-- 0x11CB
		when 004556 => D <= "01010010";	-- 0x11CC
		when 004557 => D <= "01001000";	-- 0x11CD
		when 004558 => D <= "01001111";	-- 0x11CE
		when 004559 => D <= "01001100";	-- 0x11CF
		when 004560 => D <= "11000101";	-- 0x11D0
		when 004561 => D <= "10001100";	-- 0x11D1
		when 004562 => D <= "00000000";	-- 0x11D2
		when 004563 => D <= "00000010";	-- 0x11D3
		when 004564 => D <= "01010010";	-- 0x11D4
		when 004565 => D <= "01010101";	-- 0x11D5
		when 004566 => D <= "01000101";	-- 0x11D6
		when 004567 => D <= "01000011";	-- 0x11D7
		when 004568 => D <= "01001011";	-- 0x11D8
		when 004569 => D <= "01001011";	-- 0x11D9
		when 004570 => D <= "01000101";	-- 0x11DA
		when 004571 => D <= "01001000";	-- 0x11DB
		when 004572 => D <= "11010010";	-- 0x11DC
		when 004573 => D <= "10001101";	-- 0x11DD
		when 004574 => D <= "00000000";	-- 0x11DE
		when 004575 => D <= "00000010";	-- 0x11DF
		when 004576 => D <= "01010010";	-- 0x11E0
		when 004577 => D <= "01010101";	-- 0x11E1
		when 004578 => D <= "01000101";	-- 0x11E2
		when 004579 => D <= "01000011";	-- 0x11E3
		when 004580 => D <= "01001011";	-- 0x11E4
		when 004581 => D <= "01010111";	-- 0x11E5
		when 004582 => D <= "01000001";	-- 0x11E6
		when 004583 => D <= "01000101";	-- 0x11E7
		when 004584 => D <= "01010010";	-- 0x11E8
		when 004585 => D <= "01010100";	-- 0x11E9
		when 004586 => D <= "11010011";	-- 0x11EA
		when 004587 => D <= "10000001";	-- 0x11EB
		when 004588 => D <= "00000000";	-- 0x11EC
		when 004589 => D <= "00000010";	-- 0x11ED
		when 004590 => D <= "01010110";	-- 0x11EE
		when 004591 => D <= "01001111";	-- 0x11EF
		when 004592 => D <= "01010010";	-- 0x11F0
		when 004593 => D <= "01010111";	-- 0x11F1
		when 004594 => D <= "01000001";	-- 0x11F2
		when 004595 => D <= "01000101";	-- 0x11F3
		when 004596 => D <= "01010010";	-- 0x11F4
		when 004597 => D <= "01010100";	-- 0x11F5
		when 004598 => D <= "11010011";	-- 0x11F6
		when 004599 => D <= "10000010";	-- 0x11F7
		when 004600 => D <= "00000000";	-- 0x11F8
		when 004601 => D <= "00000010";	-- 0x11F9
		when 004602 => D <= "01010011";	-- 0x11FA
		when 004603 => D <= "01000011";	-- 0x11FB
		when 004604 => D <= "01001000";	-- 0x11FC
		when 004605 => D <= "01010010";	-- 0x11FD
		when 004606 => D <= "00110001";	-- 0x11FE
		when 004607 => D <= "00110110";	-- 0x11FF
		when 004608 => D <= "01010100";	-- 0x1200
		when 004609 => D <= "01000101";	-- 0x1201
		when 004610 => D <= "11001100";	-- 0x1202
		when 004611 => D <= "10011000";	-- 0x1203
		when 004612 => D <= "00000000";	-- 0x1204
		when 004613 => D <= "00000010";	-- 0x1205
		when 004614 => D <= "01001100";	-- 0x1206
		when 004615 => D <= "01001001";	-- 0x1207
		when 004616 => D <= "01001110";	-- 0x1208
		when 004617 => D <= "01001011";	-- 0x1209
		when 004618 => D <= "11010011";	-- 0x120A
		when 004619 => D <= "10000011";	-- 0x120B
		when 004620 => D <= "00000000";	-- 0x120C
		when 004621 => D <= "00000010";	-- 0x120D
		when 004622 => D <= "01010010";	-- 0x120E
		when 004623 => D <= "01000101";	-- 0x120F
		when 004624 => D <= "01000011";	-- 0x1210
		when 004625 => D <= "01001000";	-- 0x1211
		when 004626 => D <= "01010100";	-- 0x1212
		when 004627 => D <= "11010011";	-- 0x1213
		when 004628 => D <= "10000100";	-- 0x1214
		when 004629 => D <= "00000000";	-- 0x1215
		when 004630 => D <= "00000010";	-- 0x1216
		when 004631 => D <= "01010011";	-- 0x1217
		when 004632 => D <= "01010100";	-- 0x1218
		when 004633 => D <= "01001001";	-- 0x1219
		when 004634 => D <= "01000110";	-- 0x121A
		when 004635 => D <= "01010100";	-- 0x121B
		when 004636 => D <= "01000001";	-- 0x121C
		when 004637 => D <= "11000010";	-- 0x121D
		when 004638 => D <= "10000101";	-- 0x121E
		when 004639 => D <= "00000000";	-- 0x121F
		when 004640 => D <= "00000010";	-- 0x1220
		when 004641 => D <= "01010011";	-- 0x1221
		when 004642 => D <= "11000001";	-- 0x1222
		when 004643 => D <= "10000101";	-- 0x1223
		when 004644 => D <= "00000000";	-- 0x1224
		when 004645 => D <= "00000010";	-- 0x1225
		when 004646 => D <= "01010011";	-- 0x1226
		when 004647 => D <= "01010100";	-- 0x1227
		when 004648 => D <= "01001001";	-- 0x1228
		when 004649 => D <= "01000110";	-- 0x1229
		when 004650 => D <= "01010100";	-- 0x122A
		when 004651 => D <= "01001000";	-- 0x122B
		when 004652 => D <= "01001111";	-- 0x122C
		when 004653 => D <= "01000011";	-- 0x122D
		when 004654 => D <= "11001000";	-- 0x122E
		when 004655 => D <= "10000110";	-- 0x122F
		when 004656 => D <= "00000000";	-- 0x1230
		when 004657 => D <= "00000010";	-- 0x1231
		when 004658 => D <= "01010011";	-- 0x1232
		when 004659 => D <= "11001000";	-- 0x1233
		when 004660 => D <= "10000110";	-- 0x1234
		when 004661 => D <= "00000000";	-- 0x1235
		when 004662 => D <= "00000010";	-- 0x1236
		when 004663 => D <= "01010110";	-- 0x1237
		when 004664 => D <= "11001001";	-- 0x1238
		when 004665 => D <= "10000111";	-- 0x1239
		when 004666 => D <= "00000000";	-- 0x123A
		when 004667 => D <= "00000010";	-- 0x123B
		when 004668 => D <= "01011010";	-- 0x123C
		when 004669 => D <= "11001001";	-- 0x123D
		when 004670 => D <= "10001000";	-- 0x123E
		when 004671 => D <= "00000000";	-- 0x123F
		when 004672 => D <= "00000010";	-- 0x1240
		when 004673 => D <= "01000100";	-- 0x1241
		when 004674 => D <= "01010010";	-- 0x1242
		when 004675 => D <= "01010101";	-- 0x1243
		when 004676 => D <= "01000011";	-- 0x1244
		when 004677 => D <= "01001011";	-- 0x1245
		when 004678 => D <= "01000101";	-- 0x1246
		when 004679 => D <= "01011010";	-- 0x1247
		when 004680 => D <= "01000101";	-- 0x1248
		when 004681 => D <= "01001001";	-- 0x1249
		when 004682 => D <= "01001100";	-- 0x124A
		when 004683 => D <= "11000101";	-- 0x124B
		when 004684 => D <= "10001110";	-- 0x124C
		when 004685 => D <= "00000000";	-- 0x124D
		when 004686 => D <= "00000010";	-- 0x124E
		when 004687 => D <= "01000100";	-- 0x124F
		when 004688 => D <= "11011010";	-- 0x1250
		when 004689 => D <= "10001110";	-- 0x1251
		when 004690 => D <= "00000000";	-- 0x1252
		when 004691 => D <= "00000010";	-- 0x1253
		when 004692 => D <= "01001101";	-- 0x1254
		when 004693 => D <= "01001001";	-- 0x1255
		when 004694 => D <= "01010100";	-- 0x1256
		when 004695 => D <= "01010100";	-- 0x1257
		when 004696 => D <= "11000101";	-- 0x1258
		when 004697 => D <= "10001111";	-- 0x1259
		when 004698 => D <= "00000000";	-- 0x125A
		when 004699 => D <= "00000010";	-- 0x125B
		when 004700 => D <= "01000001";	-- 0x125C
		when 004701 => D <= "01010101";	-- 0x125D
		when 004702 => D <= "01000110";	-- 0x125E
		when 004703 => D <= "01011000";	-- 0x125F
		when 004704 => D <= "11011001";	-- 0x1260
		when 004705 => D <= "10010000";	-- 0x1261
		when 004706 => D <= "00000000";	-- 0x1262
		when 004707 => D <= "00000010";	-- 0x1263
		when 004708 => D <= "01000001";	-- 0x1264
		when 004709 => D <= "01010101";	-- 0x1265
		when 004710 => D <= "01000110";	-- 0x1266
		when 004711 => D <= "01001011";	-- 0x1267
		when 004712 => D <= "01010101";	-- 0x1268
		when 004713 => D <= "01010010";	-- 0x1269
		when 004714 => D <= "11010011";	-- 0x126A
		when 004715 => D <= "10010001";	-- 0x126B
		when 004716 => D <= "00000000";	-- 0x126C
		when 004717 => D <= "00000010";	-- 0x126D
		when 004718 => D <= "01000001";	-- 0x126E
		when 004719 => D <= "11001011";	-- 0x126F
		when 004720 => D <= "10010001";	-- 0x1270
		when 004721 => D <= "00000000";	-- 0x1271
		when 004722 => D <= "00000010";	-- 0x1272
		when 004723 => D <= "01001100";	-- 0x1273
		when 004724 => D <= "01001111";	-- 0x1274
		when 004725 => D <= "01000101";	-- 0x1275
		when 004726 => D <= "01010011";	-- 0x1276
		when 004727 => D <= "01000011";	-- 0x1277
		when 004728 => D <= "01001000";	-- 0x1278
		when 004729 => D <= "01000101";	-- 0x1279
		when 004730 => D <= "01000010";	-- 0x127A
		when 004731 => D <= "01001001";	-- 0x127B
		when 004732 => D <= "01001100";	-- 0x127C
		when 004733 => D <= "11000100";	-- 0x127D
		when 004734 => D <= "10010010";	-- 0x127E
		when 004735 => D <= "00000000";	-- 0x127F
		when 004736 => D <= "00000010";	-- 0x1280
		when 004737 => D <= "01001100";	-- 0x1281
		when 004738 => D <= "11000010";	-- 0x1282
		when 004739 => D <= "10010010";	-- 0x1283
		when 004740 => D <= "00000000";	-- 0x1284
		when 004741 => D <= "00000010";	-- 0x1285
		when 004742 => D <= "01000010";	-- 0x1286
		when 004743 => D <= "01001100";	-- 0x1287
		when 004744 => D <= "01001001";	-- 0x1288
		when 004745 => D <= "01001110";	-- 0x1289
		when 004746 => D <= "01001011";	-- 0x128A
		when 004747 => D <= "01000101";	-- 0x128B
		when 004748 => D <= "11010010";	-- 0x128C
		when 004749 => D <= "10010111";	-- 0x128D
		when 004750 => D <= "00000000";	-- 0x128E
		when 004751 => D <= "00000010";	-- 0x128F
		when 004752 => D <= "01000100";	-- 0x1290
		when 004753 => D <= "01010010";	-- 0x1291
		when 004754 => D <= "01010101";	-- 0x1292
		when 004755 => D <= "01000011";	-- 0x1293
		when 004756 => D <= "01001011";	-- 0x1294
		when 004757 => D <= "11000101";	-- 0x1295
		when 004758 => D <= "10011001";	-- 0x1296
		when 004759 => D <= "00000000";	-- 0x1297
		when 004760 => D <= "00000010";	-- 0x1298
		when 004761 => D <= "01000100";	-- 0x1299
		when 004762 => D <= "11010010";	-- 0x129A
		when 004763 => D <= "10011001";	-- 0x129B
		when 004764 => D <= "00000000";	-- 0x129C
		when 004765 => D <= "00000010";	-- 0x129D
		when 004766 => D <= "01011010";	-- 0x129E
		when 004767 => D <= "01000101";	-- 0x129F
		when 004768 => D <= "01001001";	-- 0x12A0
		when 004769 => D <= "01000011";	-- 0x12A1
		when 004770 => D <= "01001000";	-- 0x12A2
		when 004771 => D <= "01000101";	-- 0x12A3
		when 004772 => D <= "11001110";	-- 0x12A4
		when 004773 => D <= "10011010";	-- 0x12A5
		when 004774 => D <= "00000000";	-- 0x12A6
		when 004775 => D <= "00000010";	-- 0x12A7
		when 004776 => D <= "01001100";	-- 0x12A8
		when 004777 => D <= "01001001";	-- 0x12A9
		when 004778 => D <= "01001110";	-- 0x12AA
		when 004779 => D <= "01001001";	-- 0x12AB
		when 004780 => D <= "11000101";	-- 0x12AC
		when 004781 => D <= "10011100";	-- 0x12AD
		when 004782 => D <= "00000000";	-- 0x12AE
		when 004783 => D <= "00000010";	-- 0x12AF
		when 004784 => D <= "01010011";	-- 0x12B0
		when 004785 => D <= "01000101";	-- 0x12B1
		when 004786 => D <= "01001001";	-- 0x12B2
		when 004787 => D <= "01010100";	-- 0x12B3
		when 004788 => D <= "11000101";	-- 0x12B4
		when 004789 => D <= "10011101";	-- 0x12B5
		when 004790 => D <= "00000000";	-- 0x12B6
		when 004791 => D <= "00000010";	-- 0x12B7
		when 004792 => D <= "01010000";	-- 0x12B8
		when 004793 => D <= "01010010";	-- 0x12B9
		when 004794 => D <= "01010101";	-- 0x12BA
		when 004795 => D <= "01000101";	-- 0x12BB
		when 004796 => D <= "01000110";	-- 0x12BC
		when 004797 => D <= "11000101";	-- 0x12BD
		when 004798 => D <= "10011110";	-- 0x12BE
		when 004799 => D <= "00000000";	-- 0x12BF
		when 004800 => D <= "00000010";	-- 0x12C0
		when 004801 => D <= "01010111";	-- 0x12C1
		when 004802 => D <= "01000101";	-- 0x12C2
		when 004803 => D <= "01001110";	-- 0x12C3
		when 004804 => D <= "01001110";	-- 0x12C4
		when 004805 => D <= "01010111";	-- 0x12C5
		when 004806 => D <= "01000001";	-- 0x12C6
		when 004807 => D <= "01001000";	-- 0x12C7
		when 004808 => D <= "11010010";	-- 0x12C8
		when 004809 => D <= "10011111";	-- 0x12C9
		when 004810 => D <= "00000000";	-- 0x12CA
		when 004811 => D <= "00000010";	-- 0x12CB
		when 004812 => D <= "01010111";	-- 0x12CC
		when 004813 => D <= "11010111";	-- 0x12CD
		when 004814 => D <= "10011111";	-- 0x12CE
		when 004815 => D <= "00000000";	-- 0x12CF
		when 004816 => D <= "00000010";	-- 0x12D0
		when 004817 => D <= "01010111";	-- 0x12D1
		when 004818 => D <= "01000101";	-- 0x12D2
		when 004819 => D <= "01001110";	-- 0x12D3
		when 004820 => D <= "01001110";	-- 0x12D4
		when 004821 => D <= "01000110";	-- 0x12D5
		when 004822 => D <= "01000001";	-- 0x12D6
		when 004823 => D <= "01001100";	-- 0x12D7
		when 004824 => D <= "01010011";	-- 0x12D8
		when 004825 => D <= "01000011";	-- 0x12D9
		when 004826 => D <= "11001000";	-- 0x12DA
		when 004827 => D <= "10100000";	-- 0x12DB
		when 004828 => D <= "00000000";	-- 0x12DC
		when 004829 => D <= "00000010";	-- 0x12DD
		when 004830 => D <= "01010111";	-- 0x12DE
		when 004831 => D <= "11000110";	-- 0x12DF
		when 004832 => D <= "10100000";	-- 0x12E0
		when 004833 => D <= "00000000";	-- 0x12E1
		when 004834 => D <= "00000010";	-- 0x12E2
		when 004835 => D <= "01010011";	-- 0x12E3
		when 004836 => D <= "01001111";	-- 0x12E4
		when 004837 => D <= "01001100";	-- 0x12E5
		when 004838 => D <= "01000001";	-- 0x12E6
		when 004839 => D <= "01001110";	-- 0x12E7
		when 004840 => D <= "01000111";	-- 0x12E8
		when 004841 => D <= "11000101";	-- 0x12E9
		when 004842 => D <= "10100100";	-- 0x12EA
		when 004843 => D <= "00000000";	-- 0x12EB
		when 004844 => D <= "00000010";	-- 0x12EC
		when 004845 => D <= "01000100";	-- 0x12ED
		when 004846 => D <= "01010010";	-- 0x12EE
		when 004847 => D <= "01010101";	-- 0x12EF
		when 004848 => D <= "01000011";	-- 0x12F0
		when 004849 => D <= "01001011";	-- 0x12F1
		when 004850 => D <= "01000001";	-- 0x12F2
		when 004851 => D <= "11001110";	-- 0x12F3
		when 004852 => D <= "10100010";	-- 0x12F4
		when 004853 => D <= "00000000";	-- 0x12F5
		when 004854 => D <= "00000010";	-- 0x12F6
		when 004855 => D <= "01000100";	-- 0x12F7
		when 004856 => D <= "01010010";	-- 0x12F8
		when 004857 => D <= "01010101";	-- 0x12F9
		when 004858 => D <= "01000011";	-- 0x12FA
		when 004859 => D <= "01001011";	-- 0x12FB
		when 004860 => D <= "01000001";	-- 0x12FC
		when 004861 => D <= "01010101";	-- 0x12FD
		when 004862 => D <= "11010011";	-- 0x12FE
		when 004863 => D <= "10100011";	-- 0x12FF
		when 004864 => D <= "00000000";	-- 0x1300
		when 004865 => D <= "00000010";	-- 0x1301
		when 004866 => D <= "01000010";	-- 0x1302
		when 004867 => D <= "01001001";	-- 0x1303
		when 004868 => D <= "01001100";	-- 0x1304
		when 004869 => D <= "11000100";	-- 0x1305
		when 004870 => D <= "10100101";	-- 0x1306
		when 004871 => D <= "00000000";	-- 0x1307
		when 004872 => D <= "00000010";	-- 0x1308
		when 004873 => D <= "01001100";	-- 0x1309
		when 004874 => D <= "01001111";	-- 0x130A
		when 004875 => D <= "01000101";	-- 0x130B
		when 004876 => D <= "01010011";	-- 0x130C
		when 004877 => D <= "01000011";	-- 0x130D
		when 004878 => D <= "01001000";	-- 0x130E
		when 004879 => D <= "01000101";	-- 0x130F
		when 004880 => D <= "01010011";	-- 0x1310
		when 004881 => D <= "01000011";	-- 0x1311
		when 004882 => D <= "01001000";	-- 0x1312
		when 004883 => D <= "01001001";	-- 0x1313
		when 004884 => D <= "01010010";	-- 0x1314
		when 004885 => D <= "11001101";	-- 0x1315
		when 004886 => D <= "10100110";	-- 0x1316
		when 004887 => D <= "00000000";	-- 0x1317
		when 004888 => D <= "00000010";	-- 0x1318
		when 004889 => D <= "01001100";	-- 0x1319
		when 004890 => D <= "11010011";	-- 0x131A
		when 004891 => D <= "10100110";	-- 0x131B
		when 004892 => D <= "00000000";	-- 0x131C
		when 004893 => D <= "00000010";	-- 0x131D
		when 004894 => D <= "01000001";	-- 0x131E
		when 004895 => D <= "01010101";	-- 0x131F
		when 004896 => D <= "01000110";	-- 0x1320
		when 004897 => D <= "11011000";	-- 0x1321
		when 004898 => D <= "10100111";	-- 0x1322
		when 004899 => D <= "00000000";	-- 0x1323
		when 004900 => D <= "00000010";	-- 0x1324
		when 004901 => D <= "01000001";	-- 0x1325
		when 004902 => D <= "01010101";	-- 0x1326
		when 004903 => D <= "01000110";	-- 0x1327
		when 004904 => D <= "11011001";	-- 0x1328
		when 004905 => D <= "10101000";	-- 0x1329
		when 004906 => D <= "00000000";	-- 0x132A
		when 004907 => D <= "00000010";	-- 0x132B
		when 004908 => D <= "01001100";	-- 0x132C
		when 004909 => D <= "01000101";	-- 0x132D
		when 004910 => D <= "01010010";	-- 0x132E
		when 004911 => D <= "01001110";	-- 0x132F
		when 004912 => D <= "11000101";	-- 0x1330
		when 004913 => D <= "10001001";	-- 0x1331
		when 004914 => D <= "00000000";	-- 0x1332
		when 004915 => D <= "00000010";	-- 0x1333
		when 004916 => D <= "01000110";	-- 0x1334
		when 004917 => D <= "01001100";	-- 0x1335
		when 004918 => D <= "01001001";	-- 0x1336
		when 004919 => D <= "11010000";	-- 0x1337
		when 004920 => D <= "10101001";	-- 0x1338
		when 004921 => D <= "00000000";	-- 0x1339
		when 004922 => D <= "00000010";	-- 0x133A
		when 004923 => D <= "01001101";	-- 0x133B
		when 004924 => D <= "01000101";	-- 0x133C
		when 004925 => D <= "11001101";	-- 0x133D
		when 004926 => D <= "10101010";	-- 0x133E
		when 004927 => D <= "00000000";	-- 0x133F
		when 004928 => D <= "00000010";	-- 0x1340
		when 004929 => D <= "01010011";	-- 0x1341
		when 004930 => D <= "01010100";	-- 0x1342
		when 004931 => D <= "01001001";	-- 0x1343
		when 004932 => D <= "01000110";	-- 0x1344
		when 004933 => D <= "11010100";	-- 0x1345
		when 004934 => D <= "10101011";	-- 0x1346
		when 004935 => D <= "00000000";	-- 0x1347
		when 004936 => D <= "00000010";	-- 0x1348
		when 004937 => D <= "01010100";	-- 0x1349
		when 004938 => D <= "01000101";	-- 0x134A
		when 004939 => D <= "01010011";	-- 0x134B
		when 004940 => D <= "11010100";	-- 0x134C
		when 004941 => D <= "10101100";	-- 0x134D
		when 004942 => D <= "00000000";	-- 0x134E
		when 004943 => D <= "00000010";	-- 0x134F
		when 004944 => D <= "01010110";	-- 0x1350
		when 004945 => D <= "01000101";	-- 0x1351
		when 004946 => D <= "01010010";	-- 0x1352
		when 004947 => D <= "01000111";	-- 0x1353
		when 004948 => D <= "01001001";	-- 0x1354
		when 004949 => D <= "01010011";	-- 0x1355
		when 004950 => D <= "11010011";	-- 0x1356
		when 004951 => D <= "10100001";	-- 0x1357
		when 004952 => D <= "00000000";	-- 0x1358
		when 004953 => D <= "00000010";	-- 0x1359
		when 004954 => D <= "01001100";	-- 0x135A
		when 004955 => D <= "01000001";	-- 0x135B
		when 004956 => D <= "01000100";	-- 0x135C
		when 004957 => D <= "11000101";	-- 0x135D
		when 004958 => D <= "10010011";	-- 0x135E
		when 004959 => D <= "00000000";	-- 0x135F
		when 004960 => D <= "00000010";	-- 0x1360
		when 004961 => D <= "01011010";	-- 0x1361
		when 004962 => D <= "01000101";	-- 0x1362
		when 004963 => D <= "01001001";	-- 0x1363
		when 004964 => D <= "01000111";	-- 0x1364
		when 004965 => D <= "11000101";	-- 0x1365
		when 004966 => D <= "10010100";	-- 0x1366
		when 004967 => D <= "00000000";	-- 0x1367
		when 004968 => D <= "00000010";	-- 0x1368
		when 004969 => D <= "01000010";	-- 0x1369
		when 004970 => D <= "01000101";	-- 0x136A
		when 004971 => D <= "01010111";	-- 0x136B
		when 004972 => D <= "01000001";	-- 0x136C
		when 004973 => D <= "01001000";	-- 0x136D
		when 004974 => D <= "01010010";	-- 0x136E
		when 004975 => D <= "11000101";	-- 0x136F
		when 004976 => D <= "10010101";	-- 0x1370
		when 004977 => D <= "00000000";	-- 0x1371
		when 004978 => D <= "00000010";	-- 0x1372
		when 004979 => D <= "01000011";	-- 0x1373
		when 004980 => D <= "01000001";	-- 0x1374
		when 004981 => D <= "01001100";	-- 0x1375
		when 004982 => D <= "11001100";	-- 0x1376
		when 004983 => D <= "10101101";	-- 0x1377
		when 004984 => D <= "00000000";	-- 0x1378
		when 004985 => D <= "00000010";	-- 0x1379
		when 004986 => D <= "01000011";	-- 0x137A
		when 004987 => D <= "01001100";	-- 0x137B
		when 004988 => D <= "01010010";	-- 0x137C
		when 004989 => D <= "01001001";	-- 0x137D
		when 004990 => D <= "01001110";	-- 0x137E
		when 004991 => D <= "11010110";	-- 0x137F
		when 004992 => D <= "10101110";	-- 0x1380
		when 004993 => D <= "00000000";	-- 0x1381
		when 004994 => D <= "00000010";	-- 0x1382
		when 004995 => D <= "00000000";	-- 0x1383
		when 004996 => D <= "00000000";	-- 0x1384
		when 004997 => D <= "11001101";	-- 0x1385
		when 004998 => D <= "00100010";	-- 0x1386
		when 004999 => D <= "00111100";	-- 0x1387
		when 005000 => D <= "11011010";	-- 0x1388
		when 005001 => D <= "01101110";	-- 0x1389
		when 005002 => D <= "00111111";	-- 0x138A
		when 005003 => D <= "11001101";	-- 0x138B
		when 005004 => D <= "11111010";	-- 0x138C
		when 005005 => D <= "00100010";	-- 0x138D
		when 005006 => D <= "11001101";	-- 0x138E
		when 005007 => D <= "01011110";	-- 0x138F
		when 005008 => D <= "00100100";	-- 0x1390
		when 005009 => D <= "11001001";	-- 0x1391
		when 005010 => D <= "11001101";	-- 0x1392
		when 005011 => D <= "00100010";	-- 0x1393
		when 005012 => D <= "00111100";	-- 0x1394
		when 005013 => D <= "11011010";	-- 0x1395
		when 005014 => D <= "01101110";	-- 0x1396
		when 005015 => D <= "00111111";	-- 0x1397
		when 005016 => D <= "11001101";	-- 0x1398
		when 005017 => D <= "01011110";	-- 0x1399
		when 005018 => D <= "00100100";	-- 0x139A
		when 005019 => D <= "11001001";	-- 0x139B
		when 005020 => D <= "11001101";	-- 0x139C
		when 005021 => D <= "00100010";	-- 0x139D
		when 005022 => D <= "00111100";	-- 0x139E
		when 005023 => D <= "11011010";	-- 0x139F
		when 005024 => D <= "01101110";	-- 0x13A0
		when 005025 => D <= "00111111";	-- 0x13A1
		when 005026 => D <= "11001101";	-- 0x13A2
		when 005027 => D <= "01100001";	-- 0x13A3
		when 005028 => D <= "00100100";	-- 0x13A4
		when 005029 => D <= "11001001";	-- 0x13A5
		when 005030 => D <= "11001101";	-- 0x13A6
		when 005031 => D <= "00100010";	-- 0x13A7
		when 005032 => D <= "00111100";	-- 0x13A8
		when 005033 => D <= "11011010";	-- 0x13A9
		when 005034 => D <= "01101110";	-- 0x13AA
		when 005035 => D <= "00111111";	-- 0x13AB
		when 005036 => D <= "11001101";	-- 0x13AC
		when 005037 => D <= "10101111";	-- 0x13AD
		when 005038 => D <= "00100100";	-- 0x13AE
		when 005039 => D <= "11001001";	-- 0x13AF
		when 005040 => D <= "11001101";	-- 0x13B0
		when 005041 => D <= "00100010";	-- 0x13B1
		when 005042 => D <= "00111100";	-- 0x13B2
		when 005043 => D <= "11011010";	-- 0x13B3
		when 005044 => D <= "01101110";	-- 0x13B4
		when 005045 => D <= "00111111";	-- 0x13B5
		when 005046 => D <= "11001101";	-- 0x13B6
		when 005047 => D <= "11111010";	-- 0x13B7
		when 005048 => D <= "00100010";	-- 0x13B8
		when 005049 => D <= "11001101";	-- 0x13B9
		when 005050 => D <= "10101111";	-- 0x13BA
		when 005051 => D <= "00100100";	-- 0x13BB
		when 005052 => D <= "11001001";	-- 0x13BC
		when 005053 => D <= "11001101";	-- 0x13BD
		when 005054 => D <= "00100010";	-- 0x13BE
		when 005055 => D <= "00111100";	-- 0x13BF
		when 005056 => D <= "11011010";	-- 0x13C0
		when 005057 => D <= "01101110";	-- 0x13C1
		when 005058 => D <= "00111111";	-- 0x13C2
		when 005059 => D <= "11100101";	-- 0x13C3
		when 005060 => D <= "11001101";	-- 0x13C4
		when 005061 => D <= "00100010";	-- 0x13C5
		when 005062 => D <= "00111100";	-- 0x13C6
		when 005063 => D <= "11010001";	-- 0x13C7
		when 005064 => D <= "11101011";	-- 0x13C8
		when 005065 => D <= "11011010";	-- 0x13C9
		when 005066 => D <= "01101110";	-- 0x13CA
		when 005067 => D <= "00111111";	-- 0x13CB
		when 005068 => D <= "11001101";	-- 0x13CC
		when 005069 => D <= "01111010";	-- 0x13CD
		when 005070 => D <= "00100001";	-- 0x13CE
		when 005071 => D <= "11001101";	-- 0x13CF
		when 005072 => D <= "00100010";	-- 0x13D0
		when 005073 => D <= "00111100";	-- 0x13D1
		when 005074 => D <= "11011010";	-- 0x13D2
		when 005075 => D <= "01101110";	-- 0x13D3
		when 005076 => D <= "00111111";	-- 0x13D4
		when 005077 => D <= "11100101";	-- 0x13D5
		when 005078 => D <= "11001101";	-- 0x13D6
		when 005079 => D <= "00100010";	-- 0x13D7
		when 005080 => D <= "00111100";	-- 0x13D8
		when 005081 => D <= "11010001";	-- 0x13D9
		when 005082 => D <= "11101011";	-- 0x13DA
		when 005083 => D <= "11011010";	-- 0x13DB
		when 005084 => D <= "01101110";	-- 0x13DC
		when 005085 => D <= "00111111";	-- 0x13DD
		when 005086 => D <= "11001101";	-- 0x13DE
		when 005087 => D <= "10001010";	-- 0x13DF
		when 005088 => D <= "00100001";	-- 0x13E0
		when 005089 => D <= "11001001";	-- 0x13E1
		when 005090 => D <= "11001101";	-- 0x13E2
		when 005091 => D <= "00100010";	-- 0x13E3
		when 005092 => D <= "00111100";	-- 0x13E4
		when 005093 => D <= "11011010";	-- 0x13E5
		when 005094 => D <= "01101110";	-- 0x13E6
		when 005095 => D <= "00111111";	-- 0x13E7
		when 005096 => D <= "01111101";	-- 0x13E8
		when 005097 => D <= "00110010";	-- 0x13E9
		when 005098 => D <= "01000111";	-- 0x13EA
		when 005099 => D <= "10000000";	-- 0x13EB
		when 005100 => D <= "00110010";	-- 0x13EC
		when 005101 => D <= "01000110";	-- 0x13ED
		when 005102 => D <= "10000000";	-- 0x13EE
		when 005103 => D <= "11001101";	-- 0x13EF
		when 005104 => D <= "00100010";	-- 0x13F0
		when 005105 => D <= "00111100";	-- 0x13F1
		when 005106 => D <= "11011010";	-- 0x13F2
		when 005107 => D <= "01101110";	-- 0x13F3
		when 005108 => D <= "00111111";	-- 0x13F4
		when 005109 => D <= "01111101";	-- 0x13F5
		when 005110 => D <= "00110010";	-- 0x13F6
		when 005111 => D <= "01000101";	-- 0x13F7
		when 005112 => D <= "10000000";	-- 0x13F8
		when 005113 => D <= "11001101";	-- 0x13F9
		when 005114 => D <= "01011000";	-- 0x13FA
		when 005115 => D <= "00100001";	-- 0x13FB
		when 005116 => D <= "11001001";	-- 0x13FC
		when 005117 => D <= "11001101";	-- 0x13FD
		when 005118 => D <= "11010010";	-- 0x13FE
		when 005119 => D <= "00100100";	-- 0x13FF
		when 005120 => D <= "11001001";	-- 0x1400
		when 005121 => D <= "11001101";	-- 0x1401
		when 005122 => D <= "11001011";	-- 0x1402
		when 005123 => D <= "00100100";	-- 0x1403
		when 005124 => D <= "11001001";	-- 0x1404
		when 005125 => D <= "11001101";	-- 0x1405
		when 005126 => D <= "11011010";	-- 0x1406
		when 005127 => D <= "00100100";	-- 0x1407
		when 005128 => D <= "11001001";	-- 0x1408
		when 005129 => D <= "11001101";	-- 0x1409
		when 005130 => D <= "11110110";	-- 0x140A
		when 005131 => D <= "00100100";	-- 0x140B
		when 005132 => D <= "11001001";	-- 0x140C
		when 005133 => D <= "00101010";	-- 0x140D
		when 005134 => D <= "01000011";	-- 0x140E
		when 005135 => D <= "10000011";	-- 0x140F
		when 005136 => D <= "11011101";	-- 0x1410
		when 005137 => D <= "01111110";	-- 0x1411
		when 005138 => D <= "00000000";	-- 0x1412
		when 005139 => D <= "01110111";	-- 0x1413
		when 005140 => D <= "10110111";	-- 0x1414
		when 005141 => D <= "00101000";	-- 0x1415
		when 005142 => D <= "00000101";	-- 0x1416
		when 005143 => D <= "00100011";	-- 0x1417
		when 005144 => D <= "11011101";	-- 0x1418
		when 005145 => D <= "00100011";	-- 0x1419
		when 005146 => D <= "00011000";	-- 0x141A
		when 005147 => D <= "11110100";	-- 0x141B
		when 005148 => D <= "00100011";	-- 0x141C
		when 005149 => D <= "00110110";	-- 0x141D
		when 005150 => D <= "00000000";	-- 0x141E
		when 005151 => D <= "00100010";	-- 0x141F
		when 005152 => D <= "01000011";	-- 0x1420
		when 005153 => D <= "10000011";	-- 0x1421
		when 005154 => D <= "11001001";	-- 0x1422
		when 005155 => D <= "00100010";	-- 0x1423
		when 005156 => D <= "00000101";	-- 0x1424
		when 005157 => D <= "10000000";	-- 0x1425
		when 005158 => D <= "11100101";	-- 0x1426
		when 005159 => D <= "11011101";	-- 0x1427
		when 005160 => D <= "11100001";	-- 0x1428
		when 005161 => D <= "11011101";	-- 0x1429
		when 005162 => D <= "11100101";	-- 0x142A
		when 005163 => D <= "11111101";	-- 0x142B
		when 005164 => D <= "00100001";	-- 0x142C
		when 005165 => D <= "10000111";	-- 0x142D
		when 005166 => D <= "00110001";	-- 0x142E
		when 005167 => D <= "11001101";	-- 0x142F
		when 005168 => D <= "00110101";	-- 0x1430
		when 005169 => D <= "00101010";	-- 0x1431
		when 005170 => D <= "11010010";	-- 0x1432
		when 005171 => D <= "00110111";	-- 0x1433
		when 005172 => D <= "00110100";	-- 0x1434
		when 005173 => D <= "00101110";	-- 0x1435
		when 005174 => D <= "00000000";	-- 0x1436
		when 005175 => D <= "11011101";	-- 0x1437
		when 005176 => D <= "11100001";	-- 0x1438
		when 005177 => D <= "11011101";	-- 0x1439
		when 005178 => D <= "01111110";	-- 0x143A
		when 005179 => D <= "00000000";	-- 0x143B
		when 005180 => D <= "11011101";	-- 0x143C
		when 005181 => D <= "00100011";	-- 0x143D
		when 005182 => D <= "10110111";	-- 0x143E
		when 005183 => D <= "11000010";	-- 0x143F
		when 005184 => D <= "00111001";	-- 0x1440
		when 005185 => D <= "00110100";	-- 0x1441
		when 005186 => D <= "01111101";	-- 0x1442
		when 005187 => D <= "11111110";	-- 0x1443
		when 005188 => D <= "10001010";	-- 0x1444
		when 005189 => D <= "11000010";	-- 0x1445
		when 005190 => D <= "00101001";	-- 0x1446
		when 005191 => D <= "00110100";	-- 0x1447
		when 005192 => D <= "11011101";	-- 0x1448
		when 005193 => D <= "00100010";	-- 0x1449
		when 005194 => D <= "00000111";	-- 0x144A
		when 005195 => D <= "10000000";	-- 0x144B
		when 005196 => D <= "11101101";	-- 0x144C
		when 005197 => D <= "01011011";	-- 0x144D
		when 005198 => D <= "00000101";	-- 0x144E
		when 005199 => D <= "10000000";	-- 0x144F
		when 005200 => D <= "10101111";	-- 0x1450
		when 005201 => D <= "11011101";	-- 0x1451
		when 005202 => D <= "11100101";	-- 0x1452
		when 005203 => D <= "11100001";	-- 0x1453
		when 005204 => D <= "11101101";	-- 0x1454
		when 005205 => D <= "01010010";	-- 0x1455
		when 005206 => D <= "00100010";	-- 0x1456
		when 005207 => D <= "00001001";	-- 0x1457
		when 005208 => D <= "10000000";	-- 0x1458
		when 005209 => D <= "00101010";	-- 0x1459
		when 005210 => D <= "01000011";	-- 0x145A
		when 005211 => D <= "10000011";	-- 0x145B
		when 005212 => D <= "11101101";	-- 0x145C
		when 005213 => D <= "01011011";	-- 0x145D
		when 005214 => D <= "00000111";	-- 0x145E
		when 005215 => D <= "10000000";	-- 0x145F
		when 005216 => D <= "10101111";	-- 0x1460
		when 005217 => D <= "11101101";	-- 0x1461
		when 005218 => D <= "01010010";	-- 0x1462
		when 005219 => D <= "00100011";	-- 0x1463
		when 005220 => D <= "01000100";	-- 0x1464
		when 005221 => D <= "01001101";	-- 0x1465
		when 005222 => D <= "11101101";	-- 0x1466
		when 005223 => D <= "01011011";	-- 0x1467
		when 005224 => D <= "00000101";	-- 0x1468
		when 005225 => D <= "10000000";	-- 0x1469
		when 005226 => D <= "00101010";	-- 0x146A
		when 005227 => D <= "00000111";	-- 0x146B
		when 005228 => D <= "10000000";	-- 0x146C
		when 005229 => D <= "11101101";	-- 0x146D
		when 005230 => D <= "10110000";	-- 0x146E
		when 005231 => D <= "11111101";	-- 0x146F
		when 005232 => D <= "00100001";	-- 0x1470
		when 005233 => D <= "01001111";	-- 0x1471
		when 005234 => D <= "10000011";	-- 0x1472
		when 005235 => D <= "11100101";	-- 0x1473
		when 005236 => D <= "00100001";	-- 0x1474
		when 005237 => D <= "10111010";	-- 0x1475
		when 005238 => D <= "00110100";	-- 0x1476
		when 005239 => D <= "11100011";	-- 0x1477
		when 005240 => D <= "11111101";	-- 0x1478
		when 005241 => D <= "01111110";	-- 0x1479
		when 005242 => D <= "00000000";	-- 0x147A
		when 005243 => D <= "10110111";	-- 0x147B
		when 005244 => D <= "11001000";	-- 0x147C
		when 005245 => D <= "11111101";	-- 0x147D
		when 005246 => D <= "11001011";	-- 0x147E
		when 005247 => D <= "00000000";	-- 0x147F
		when 005248 => D <= "01111110";	-- 0x1480
		when 005249 => D <= "11111101";	-- 0x1481
		when 005250 => D <= "00100011";	-- 0x1482
		when 005251 => D <= "11001010";	-- 0x1483
		when 005252 => D <= "01111101";	-- 0x1484
		when 005253 => D <= "00110100";	-- 0x1485
		when 005254 => D <= "11111101";	-- 0x1486
		when 005255 => D <= "01101110";	-- 0x1487
		when 005256 => D <= "00000000";	-- 0x1488
		when 005257 => D <= "11111101";	-- 0x1489
		when 005258 => D <= "01100110";	-- 0x148A
		when 005259 => D <= "00000001";	-- 0x148B
		when 005260 => D <= "11111101";	-- 0x148C
		when 005261 => D <= "01111110";	-- 0x148D
		when 005262 => D <= "00000010";	-- 0x148E
		when 005263 => D <= "11111110";	-- 0x148F
		when 005264 => D <= "00000010";	-- 0x1490
		when 005265 => D <= "11000010";	-- 0x1491
		when 005266 => D <= "10110001";	-- 0x1492
		when 005267 => D <= "00110100";	-- 0x1493
		when 005268 => D <= "11101101";	-- 0x1494
		when 005269 => D <= "01011011";	-- 0x1495
		when 005270 => D <= "00000111";	-- 0x1496
		when 005271 => D <= "10000000";	-- 0x1497
		when 005272 => D <= "10101111";	-- 0x1498
		when 005273 => D <= "11101101";	-- 0x1499
		when 005274 => D <= "01010010";	-- 0x149A
		when 005275 => D <= "11011010";	-- 0x149B
		when 005276 => D <= "10110001";	-- 0x149C
		when 005277 => D <= "00110100";	-- 0x149D
		when 005278 => D <= "11111101";	-- 0x149E
		when 005279 => D <= "01101110";	-- 0x149F
		when 005280 => D <= "00000000";	-- 0x14A0
		when 005281 => D <= "11111101";	-- 0x14A1
		when 005282 => D <= "01100110";	-- 0x14A2
		when 005283 => D <= "00000001";	-- 0x14A3
		when 005284 => D <= "11101101";	-- 0x14A4
		when 005285 => D <= "01011011";	-- 0x14A5
		when 005286 => D <= "00001001";	-- 0x14A6
		when 005287 => D <= "10000000";	-- 0x14A7
		when 005288 => D <= "10101111";	-- 0x14A8
		when 005289 => D <= "11101101";	-- 0x14A9
		when 005290 => D <= "01010010";	-- 0x14AA
		when 005291 => D <= "11111101";	-- 0x14AB
		when 005292 => D <= "01110101";	-- 0x14AC
		when 005293 => D <= "00000000";	-- 0x14AD
		when 005294 => D <= "11111101";	-- 0x14AE
		when 005295 => D <= "01110100";	-- 0x14AF
		when 005296 => D <= "00000001";	-- 0x14B0
		when 005297 => D <= "11111101";	-- 0x14B1
		when 005298 => D <= "00100011";	-- 0x14B2
		when 005299 => D <= "11111101";	-- 0x14B3
		when 005300 => D <= "00100011";	-- 0x14B4
		when 005301 => D <= "11111101";	-- 0x14B5
		when 005302 => D <= "00100011";	-- 0x14B6
		when 005303 => D <= "11000011";	-- 0x14B7
		when 005304 => D <= "01111000";	-- 0x14B8
		when 005305 => D <= "00110100";	-- 0x14B9
		when 005306 => D <= "00101010";	-- 0x14BA
		when 005307 => D <= "01000011";	-- 0x14BB
		when 005308 => D <= "10000011";	-- 0x14BC
		when 005309 => D <= "11101101";	-- 0x14BD
		when 005310 => D <= "01011011";	-- 0x14BE
		when 005311 => D <= "00001001";	-- 0x14BF
		when 005312 => D <= "10000000";	-- 0x14C0
		when 005313 => D <= "10101111";	-- 0x14C1
		when 005314 => D <= "11101101";	-- 0x14C2
		when 005315 => D <= "01010010";	-- 0x14C3
		when 005316 => D <= "00100010";	-- 0x14C4
		when 005317 => D <= "01000011";	-- 0x14C5
		when 005318 => D <= "10000011";	-- 0x14C6
		when 005319 => D <= "11001001";	-- 0x14C7
		when 005320 => D <= "00100001";	-- 0x14C8
		when 005321 => D <= "00000000";	-- 0x14C9
		when 005322 => D <= "00000000";	-- 0x14CA
		when 005323 => D <= "00100010";	-- 0x14CB
		when 005324 => D <= "00001011";	-- 0x14CC
		when 005325 => D <= "10000000";	-- 0x14CD
		when 005326 => D <= "11001101";	-- 0x14CE
		when 005327 => D <= "11001100";	-- 0x14CF
		when 005328 => D <= "00100111";	-- 0x14D0
		when 005329 => D <= "11011101";	-- 0x14D1
		when 005330 => D <= "11100101";	-- 0x14D2
		when 005331 => D <= "00101010";	-- 0x14D3
		when 005332 => D <= "01000011";	-- 0x14D4
		when 005333 => D <= "10000011";	-- 0x14D5
		when 005334 => D <= "00100010";	-- 0x14D6
		when 005335 => D <= "00001111";	-- 0x14D7
		when 005336 => D <= "10000000";	-- 0x14D8
		when 005337 => D <= "00111110";	-- 0x14D9
		when 005338 => D <= "00000010";	-- 0x14DA
		when 005339 => D <= "11001101";	-- 0x14DB
		when 005340 => D <= "01110010";	-- 0x14DC
		when 005341 => D <= "00101011";	-- 0x14DD
		when 005342 => D <= "11010010";	-- 0x14DE
		when 005343 => D <= "00001011";	-- 0x14DF
		when 005344 => D <= "00110101";	-- 0x14E0
		when 005345 => D <= "11011101";	-- 0x14E1
		when 005346 => D <= "11100001";	-- 0x14E2
		when 005347 => D <= "11011101";	-- 0x14E3
		when 005348 => D <= "11100101";	-- 0x14E4
		when 005349 => D <= "11011101";	-- 0x14E5
		when 005350 => D <= "11100101";	-- 0x14E6
		when 005351 => D <= "11111110";	-- 0x14E7
		when 005352 => D <= "00000010";	-- 0x14E8
		when 005353 => D <= "11000010";	-- 0x14E9
		when 005354 => D <= "11101111";	-- 0x14EA
		when 005355 => D <= "00110100";	-- 0x14EB
		when 005356 => D <= "11001101";	-- 0x14EC
		when 005357 => D <= "00100011";	-- 0x14ED
		when 005358 => D <= "00110100";	-- 0x14EE
		when 005359 => D <= "11011101";	-- 0x14EF
		when 005360 => D <= "11100001";	-- 0x14F0
		when 005361 => D <= "11111101";	-- 0x14F1
		when 005362 => D <= "00100001";	-- 0x14F2
		when 005363 => D <= "01001111";	-- 0x14F3
		when 005364 => D <= "10000011";	-- 0x14F4
		when 005365 => D <= "11001101";	-- 0x14F5
		when 005366 => D <= "00110101";	-- 0x14F6
		when 005367 => D <= "00101010";	-- 0x14F7
		when 005368 => D <= "11011010";	-- 0x14F8
		when 005369 => D <= "01101110";	-- 0x14F9
		when 005370 => D <= "00111111";	-- 0x14FA
		when 005371 => D <= "00101010";	-- 0x14FB
		when 005372 => D <= "01000011";	-- 0x14FC
		when 005373 => D <= "10000011";	-- 0x14FD
		when 005374 => D <= "00100010";	-- 0x14FE
		when 005375 => D <= "00001111";	-- 0x14FF
		when 005376 => D <= "10000000";	-- 0x1500
		when 005377 => D <= "11111101";	-- 0x1501
		when 005378 => D <= "01110101";	-- 0x1502
		when 005379 => D <= "00000000";	-- 0x1503
		when 005380 => D <= "11111101";	-- 0x1504
		when 005381 => D <= "01110100";	-- 0x1505
		when 005382 => D <= "00000001";	-- 0x1506
		when 005383 => D <= "11111101";	-- 0x1507
		when 005384 => D <= "00110110";	-- 0x1508
		when 005385 => D <= "00000010";	-- 0x1509
		when 005386 => D <= "00000010";	-- 0x150A
		when 005387 => D <= "11011101";	-- 0x150B
		when 005388 => D <= "11100001";	-- 0x150C
		when 005389 => D <= "11001101";	-- 0x150D
		when 005390 => D <= "11001100";	-- 0x150E
		when 005391 => D <= "00100111";	-- 0x150F
		when 005392 => D <= "11001101";	-- 0x1510
		when 005393 => D <= "00001101";	-- 0x1511
		when 005394 => D <= "00110100";	-- 0x1512
		when 005395 => D <= "00101010";	-- 0x1513
		when 005396 => D <= "00001011";	-- 0x1514
		when 005397 => D <= "10000000";	-- 0x1515
		when 005398 => D <= "00100010";	-- 0x1516
		when 005399 => D <= "00001101";	-- 0x1517
		when 005400 => D <= "10000000";	-- 0x1518
		when 005401 => D <= "00101010";	-- 0x1519
		when 005402 => D <= "01000011";	-- 0x151A
		when 005403 => D <= "10000011";	-- 0x151B
		when 005404 => D <= "00100010";	-- 0x151C
		when 005405 => D <= "00001011";	-- 0x151D
		when 005406 => D <= "10000000";	-- 0x151E
		when 005407 => D <= "11001101";	-- 0x151F
		when 005408 => D <= "11111001";	-- 0x1520
		when 005409 => D <= "00110000";	-- 0x1521
		when 005410 => D <= "11100101";	-- 0x1522
		when 005411 => D <= "11011101";	-- 0x1523
		when 005412 => D <= "11100001";	-- 0x1524
		when 005413 => D <= "11001101";	-- 0x1525
		when 005414 => D <= "11001100";	-- 0x1526
		when 005415 => D <= "00100111";	-- 0x1527
		when 005416 => D <= "11011101";	-- 0x1528
		when 005417 => D <= "11100101";	-- 0x1529
		when 005418 => D <= "11001101";	-- 0x152A
		when 005419 => D <= "00001101";	-- 0x152B
		when 005420 => D <= "00110100";	-- 0x152C
		when 005421 => D <= "11011101";	-- 0x152D
		when 005422 => D <= "11100001";	-- 0x152E
		when 005423 => D <= "11111101";	-- 0x152F
		when 005424 => D <= "00100001";	-- 0x1530
		when 005425 => D <= "10000111";	-- 0x1531
		when 005426 => D <= "00110001";	-- 0x1532
		when 005427 => D <= "11001101";	-- 0x1533
		when 005428 => D <= "00110101";	-- 0x1534
		when 005429 => D <= "00101010";	-- 0x1535
		when 005430 => D <= "11010010";	-- 0x1536
		when 005431 => D <= "00111011";	-- 0x1537
		when 005432 => D <= "00110101";	-- 0x1538
		when 005433 => D <= "00101110";	-- 0x1539
		when 005434 => D <= "00000000";	-- 0x153A
		when 005435 => D <= "01111101";	-- 0x153B
		when 005436 => D <= "11111110";	-- 0x153C
		when 005437 => D <= "10001010";	-- 0x153D
		when 005438 => D <= "11000010";	-- 0x153E
		when 005439 => D <= "00010011";	-- 0x153F
		when 005440 => D <= "00110101";	-- 0x1540
		when 005441 => D <= "00101010";	-- 0x1541
		when 005442 => D <= "00001101";	-- 0x1542
		when 005443 => D <= "10000000";	-- 0x1543
		when 005444 => D <= "01111100";	-- 0x1544
		when 005445 => D <= "10110101";	-- 0x1545
		when 005446 => D <= "11001010";	-- 0x1546
		when 005447 => D <= "01101101";	-- 0x1547
		when 005448 => D <= "00110101";	-- 0x1548
		when 005449 => D <= "11011101";	-- 0x1549
		when 005450 => D <= "00101010";	-- 0x154A
		when 005451 => D <= "00001101";	-- 0x154B
		when 005452 => D <= "10000000";	-- 0x154C
		when 005453 => D <= "11111101";	-- 0x154D
		when 005454 => D <= "00100001";	-- 0x154E
		when 005455 => D <= "01001111";	-- 0x154F
		when 005456 => D <= "10000011";	-- 0x1550
		when 005457 => D <= "11001101";	-- 0x1551
		when 005458 => D <= "00110101";	-- 0x1552
		when 005459 => D <= "00101010";	-- 0x1553
		when 005460 => D <= "11011010";	-- 0x1554
		when 005461 => D <= "01101101";	-- 0x1555
		when 005462 => D <= "00110101";	-- 0x1556
		when 005463 => D <= "11111110";	-- 0x1557
		when 005464 => D <= "00000010";	-- 0x1558
		when 005465 => D <= "11000010";	-- 0x1559
		when 005466 => D <= "01101101";	-- 0x155A
		when 005467 => D <= "00110101";	-- 0x155B
		when 005468 => D <= "11101101";	-- 0x155C
		when 005469 => D <= "01011011";	-- 0x155D
		when 005470 => D <= "00001111";	-- 0x155E
		when 005471 => D <= "10000000";	-- 0x155F
		when 005472 => D <= "10101111";	-- 0x1560
		when 005473 => D <= "11101101";	-- 0x1561
		when 005474 => D <= "01010010";	-- 0x1562
		when 005475 => D <= "01111100";	-- 0x1563
		when 005476 => D <= "10110101";	-- 0x1564
		when 005477 => D <= "11000010";	-- 0x1565
		when 005478 => D <= "01101101";	-- 0x1566
		when 005479 => D <= "00110101";	-- 0x1567
		when 005480 => D <= "00101010";	-- 0x1568
		when 005481 => D <= "00001101";	-- 0x1569
		when 005482 => D <= "10000000";	-- 0x156A
		when 005483 => D <= "11001011";	-- 0x156B
		when 005484 => D <= "11111110";	-- 0x156C
		when 005485 => D <= "00100001";	-- 0x156D
		when 005486 => D <= "10100010";	-- 0x156E
		when 005487 => D <= "00110101";	-- 0x156F
		when 005488 => D <= "11001101";	-- 0x1570
		when 005489 => D <= "10110010";	-- 0x1571
		when 005490 => D <= "00111110";	-- 0x1572
		when 005491 => D <= "00101010";	-- 0x1573
		when 005492 => D <= "01000101";	-- 0x1574
		when 005493 => D <= "10000011";	-- 0x1575
		when 005494 => D <= "11101101";	-- 0x1576
		when 005495 => D <= "01011011";	-- 0x1577
		when 005496 => D <= "01000011";	-- 0x1578
		when 005497 => D <= "10000011";	-- 0x1579
		when 005498 => D <= "10101111";	-- 0x157A
		when 005499 => D <= "11101101";	-- 0x157B
		when 005500 => D <= "01010010";	-- 0x157C
		when 005501 => D <= "11001101";	-- 0x157D
		when 005502 => D <= "00001111";	-- 0x157E
		when 005503 => D <= "00101010";	-- 0x157F
		when 005504 => D <= "00100001";	-- 0x1580
		when 005505 => D <= "11000011";	-- 0x1581
		when 005506 => D <= "00110101";	-- 0x1582
		when 005507 => D <= "11001101";	-- 0x1583
		when 005508 => D <= "10110010";	-- 0x1584
		when 005509 => D <= "00111110";	-- 0x1585
		when 005510 => D <= "00101010";	-- 0x1586
		when 005511 => D <= "01000001";	-- 0x1587
		when 005512 => D <= "10000011";	-- 0x1588
		when 005513 => D <= "11101101";	-- 0x1589
		when 005514 => D <= "01011011";	-- 0x158A
		when 005515 => D <= "01001001";	-- 0x158B
		when 005516 => D <= "10000011";	-- 0x158C
		when 005517 => D <= "10101111";	-- 0x158D
		when 005518 => D <= "11101101";	-- 0x158E
		when 005519 => D <= "01010010";	-- 0x158F
		when 005520 => D <= "11001101";	-- 0x1590
		when 005521 => D <= "00001111";	-- 0x1591
		when 005522 => D <= "00101010";	-- 0x1592
		when 005523 => D <= "00100001";	-- 0x1593
		when 005524 => D <= "11011011";	-- 0x1594
		when 005525 => D <= "00110101";	-- 0x1595
		when 005526 => D <= "11001101";	-- 0x1596
		when 005527 => D <= "10110010";	-- 0x1597
		when 005528 => D <= "00111110";	-- 0x1598
		when 005529 => D <= "11011101";	-- 0x1599
		when 005530 => D <= "00100001";	-- 0x159A
		when 005531 => D <= "11101111";	-- 0x159B
		when 005532 => D <= "10000010";	-- 0x159C
		when 005533 => D <= "11011101";	-- 0x159D
		when 005534 => D <= "00110110";	-- 0x159E
		when 005535 => D <= "00000000";	-- 0x159F
		when 005536 => D <= "00000000";	-- 0x15A0
		when 005537 => D <= "11001001";	-- 0x15A1
		when 005538 => D <= "00001101";	-- 0x15A2
		when 005539 => D <= "00001010";	-- 0x15A3
		when 005540 => D <= "01001111";	-- 0x15A4
		when 005541 => D <= "01101011";	-- 0x15A5
		when 005542 => D <= "00100000";	-- 0x15A6
		when 005543 => D <= "01100111";	-- 0x15A7
		when 005544 => D <= "01100101";	-- 0x15A8
		when 005545 => D <= "01101100";	-- 0x15A9
		when 005546 => D <= "01100101";	-- 0x15AA
		when 005547 => D <= "01110010";	-- 0x15AB
		when 005548 => D <= "01101110";	-- 0x15AC
		when 005549 => D <= "01110100";	-- 0x15AD
		when 005550 => D <= "00101100";	-- 0x15AE
		when 005551 => D <= "00100000";	-- 0x15AF
		when 005552 => D <= "01010000";	-- 0x15B0
		when 005553 => D <= "01101100";	-- 0x15B1
		when 005554 => D <= "01100001";	-- 0x15B2
		when 005555 => D <= "01110100";	-- 0x15B3
		when 005556 => D <= "01111010";	-- 0x15B4
		when 005557 => D <= "00100000";	-- 0x15B5
		when 005558 => D <= "01111010";	-- 0x15B6
		when 005559 => D <= "01110101";	-- 0x15B7
		when 005560 => D <= "01101101";	-- 0x15B8
		when 005561 => D <= "00100000";	-- 0x15B9
		when 005562 => D <= "01101100";	-- 0x15BA
		when 005563 => D <= "01100101";	-- 0x15BB
		when 005564 => D <= "01110010";	-- 0x15BC
		when 005565 => D <= "01101110";	-- 0x15BD
		when 005566 => D <= "01100101";	-- 0x15BE
		when 005567 => D <= "01101110";	-- 0x15BF
		when 005568 => D <= "00111010";	-- 0x15C0
		when 005569 => D <= "00100000";	-- 0x15C1
		when 005570 => D <= "00000000";	-- 0x15C2
		when 005571 => D <= "00100000";	-- 0x15C3
		when 005572 => D <= "01000010";	-- 0x15C4
		when 005573 => D <= "01111001";	-- 0x15C5
		when 005574 => D <= "01110100";	-- 0x15C6
		when 005575 => D <= "01100101";	-- 0x15C7
		when 005576 => D <= "01110011";	-- 0x15C8
		when 005577 => D <= "00100000";	-- 0x15C9
		when 005578 => D <= "01110101";	-- 0x15CA
		when 005579 => D <= "01101110";	-- 0x15CB
		when 005580 => D <= "01100100";	-- 0x15CC
		when 005581 => D <= "00100000";	-- 0x15CD
		when 005582 => D <= "01100110";	-- 0x15CE
		when 005583 => D <= "01110101";	-- 0x15CF
		when 005584 => D <= "01100101";	-- 0x15D0
		when 005585 => D <= "01110010";	-- 0x15D1
		when 005586 => D <= "00100000";	-- 0x15D2
		when 005587 => D <= "01001110";	-- 0x15D3
		when 005588 => D <= "01100001";	-- 0x15D4
		when 005589 => D <= "01101101";	-- 0x15D5
		when 005590 => D <= "01100101";	-- 0x15D6
		when 005591 => D <= "01101110";	-- 0x15D7
		when 005592 => D <= "00111010";	-- 0x15D8
		when 005593 => D <= "00100000";	-- 0x15D9
		when 005594 => D <= "00000000";	-- 0x15DA
		when 005595 => D <= "00100000";	-- 0x15DB
		when 005596 => D <= "01000010";	-- 0x15DC
		when 005597 => D <= "01111001";	-- 0x15DD
		when 005598 => D <= "01110100";	-- 0x15DE
		when 005599 => D <= "01100101";	-- 0x15DF
		when 005600 => D <= "01110011";	-- 0x15E0
		when 005601 => D <= "00101110";	-- 0x15E1
		when 005602 => D <= "00001101";	-- 0x15E2
		when 005603 => D <= "00001010";	-- 0x15E3
		when 005604 => D <= "00000000";	-- 0x15E4
		when 005605 => D <= "00111010";	-- 0x15E5
		when 005606 => D <= "00000010";	-- 0x15E6
		when 005607 => D <= "10000000";	-- 0x15E7
		when 005608 => D <= "11111110";	-- 0x15E8
		when 005609 => D <= "11111111";	-- 0x15E9
		when 005610 => D <= "11000010";	-- 0x15EA
		when 005611 => D <= "11110100";	-- 0x15EB
		when 005612 => D <= "00110101";	-- 0x15EC
		when 005613 => D <= "10101111";	-- 0x15ED
		when 005614 => D <= "00110010";	-- 0x15EE
		when 005615 => D <= "00000010";	-- 0x15EF
		when 005616 => D <= "10000000";	-- 0x15F0
		when 005617 => D <= "11000011";	-- 0x15F1
		when 005618 => D <= "11110111";	-- 0x15F2
		when 005619 => D <= "00110101";	-- 0x15F3
		when 005620 => D <= "11000011";	-- 0x15F4
		when 005621 => D <= "01101110";	-- 0x15F5
		when 005622 => D <= "00111111";	-- 0x15F6
		when 005623 => D <= "11001001";	-- 0x15F7
		when 005624 => D <= "11001101";	-- 0x15F8
		when 005625 => D <= "00100010";	-- 0x15F9
		when 005626 => D <= "00111100";	-- 0x15FA
		when 005627 => D <= "11011010";	-- 0x15FB
		when 005628 => D <= "01111011";	-- 0x15FC
		when 005629 => D <= "00110110";	-- 0x15FD
		when 005630 => D <= "01111101";	-- 0x15FE
		when 005631 => D <= "10110100";	-- 0x15FF
		when 005632 => D <= "11000010";	-- 0x1600
		when 005633 => D <= "01000000";	-- 0x1601
		when 005634 => D <= "00110110";	-- 0x1602
		when 005635 => D <= "11001101";	-- 0x1603
		when 005636 => D <= "11001100";	-- 0x1604
		when 005637 => D <= "00100111";	-- 0x1605
		when 005638 => D <= "11111110";	-- 0x1606
		when 005639 => D <= "01011011";	-- 0x1607
		when 005640 => D <= "11000010";	-- 0x1608
		when 005641 => D <= "00111010";	-- 0x1609
		when 005642 => D <= "00110110";	-- 0x160A
		when 005643 => D <= "11001101";	-- 0x160B
		when 005644 => D <= "10110100";	-- 0x160C
		when 005645 => D <= "00110111";	-- 0x160D
		when 005646 => D <= "11001101";	-- 0x160E
		when 005647 => D <= "11001100";	-- 0x160F
		when 005648 => D <= "00100111";	-- 0x1610
		when 005649 => D <= "11111110";	-- 0x1611
		when 005650 => D <= "01011011";	-- 0x1612
		when 005651 => D <= "11000010";	-- 0x1613
		when 005652 => D <= "00110111";	-- 0x1614
		when 005653 => D <= "00110110";	-- 0x1615
		when 005654 => D <= "11011101";	-- 0x1616
		when 005655 => D <= "00100011";	-- 0x1617
		when 005656 => D <= "11001101";	-- 0x1618
		when 005657 => D <= "11001100";	-- 0x1619
		when 005658 => D <= "00100111";	-- 0x161A
		when 005659 => D <= "11111110";	-- 0x161B
		when 005660 => D <= "01011101";	-- 0x161C
		when 005661 => D <= "11001010";	-- 0x161D
		when 005662 => D <= "00110000";	-- 0x161E
		when 005663 => D <= "00110110";	-- 0x161F
		when 005664 => D <= "10110111";	-- 0x1620
		when 005665 => D <= "11001010";	-- 0x1621
		when 005666 => D <= "00110000";	-- 0x1622
		when 005667 => D <= "00110110";	-- 0x1623
		when 005668 => D <= "11001101";	-- 0x1624
		when 005669 => D <= "00111011";	-- 0x1625
		when 005670 => D <= "00111100";	-- 0x1626
		when 005671 => D <= "11001101";	-- 0x1627
		when 005672 => D <= "11001100";	-- 0x1628
		when 005673 => D <= "00100111";	-- 0x1629
		when 005674 => D <= "11011101";	-- 0x162A
		when 005675 => D <= "01111110";	-- 0x162B
		when 005676 => D <= "00000000";	-- 0x162C
		when 005677 => D <= "11000011";	-- 0x162D
		when 005678 => D <= "00011011";	-- 0x162E
		when 005679 => D <= "00110110";	-- 0x162F
		when 005680 => D <= "11111110";	-- 0x1630
		when 005681 => D <= "01011101";	-- 0x1631
		when 005682 => D <= "11000010";	-- 0x1632
		when 005683 => D <= "00110111";	-- 0x1633
		when 005684 => D <= "00110110";	-- 0x1634
		when 005685 => D <= "11011101";	-- 0x1635
		when 005686 => D <= "00100011";	-- 0x1636
		when 005687 => D <= "11000011";	-- 0x1637
		when 005688 => D <= "00111101";	-- 0x1638
		when 005689 => D <= "00110110";	-- 0x1639
		when 005690 => D <= "11000011";	-- 0x163A
		when 005691 => D <= "01101110";	-- 0x163B
		when 005692 => D <= "00111111";	-- 0x163C
		when 005693 => D <= "11000011";	-- 0x163D
		when 005694 => D <= "01111000";	-- 0x163E
		when 005695 => D <= "00110110";	-- 0x163F
		when 005696 => D <= "11001101";	-- 0x1640
		when 005697 => D <= "11001100";	-- 0x1641
		when 005698 => D <= "00100111";	-- 0x1642
		when 005699 => D <= "11111110";	-- 0x1643
		when 005700 => D <= "01011011";	-- 0x1644
		when 005701 => D <= "11000010";	-- 0x1645
		when 005702 => D <= "01110101";	-- 0x1646
		when 005703 => D <= "00110110";	-- 0x1647
		when 005704 => D <= "11011101";	-- 0x1648
		when 005705 => D <= "00100011";	-- 0x1649
		when 005706 => D <= "11001101";	-- 0x164A
		when 005707 => D <= "11001100";	-- 0x164B
		when 005708 => D <= "00100111";	-- 0x164C
		when 005709 => D <= "11011101";	-- 0x164D
		when 005710 => D <= "01111110";	-- 0x164E
		when 005711 => D <= "00000000";	-- 0x164F
		when 005712 => D <= "11111110";	-- 0x1650
		when 005713 => D <= "01011101";	-- 0x1651
		when 005714 => D <= "11001010";	-- 0x1652
		when 005715 => D <= "01100101";	-- 0x1653
		when 005716 => D <= "00110110";	-- 0x1654
		when 005717 => D <= "10110111";	-- 0x1655
		when 005718 => D <= "11001010";	-- 0x1656
		when 005719 => D <= "01100101";	-- 0x1657
		when 005720 => D <= "00110110";	-- 0x1658
		when 005721 => D <= "11001101";	-- 0x1659
		when 005722 => D <= "00111011";	-- 0x165A
		when 005723 => D <= "00111100";	-- 0x165B
		when 005724 => D <= "11001101";	-- 0x165C
		when 005725 => D <= "11001100";	-- 0x165D
		when 005726 => D <= "00100111";	-- 0x165E
		when 005727 => D <= "11011101";	-- 0x165F
		when 005728 => D <= "01111110";	-- 0x1660
		when 005729 => D <= "00000000";	-- 0x1661
		when 005730 => D <= "11000011";	-- 0x1662
		when 005731 => D <= "01010000";	-- 0x1663
		when 005732 => D <= "00110110";	-- 0x1664
		when 005733 => D <= "11111110";	-- 0x1665
		when 005734 => D <= "01011101";	-- 0x1666
		when 005735 => D <= "11000010";	-- 0x1667
		when 005736 => D <= "01101100";	-- 0x1668
		when 005737 => D <= "00110110";	-- 0x1669
		when 005738 => D <= "11011101";	-- 0x166A
		when 005739 => D <= "00100011";	-- 0x166B
		when 005740 => D <= "11001101";	-- 0x166C
		when 005741 => D <= "11001100";	-- 0x166D
		when 005742 => D <= "00100111";	-- 0x166E
		when 005743 => D <= "11001101";	-- 0x166F
		when 005744 => D <= "10110100";	-- 0x1670
		when 005745 => D <= "00110111";	-- 0x1671
		when 005746 => D <= "11000011";	-- 0x1672
		when 005747 => D <= "01111000";	-- 0x1673
		when 005748 => D <= "00110110";	-- 0x1674
		when 005749 => D <= "11000011";	-- 0x1675
		when 005750 => D <= "01101110";	-- 0x1676
		when 005751 => D <= "00111111";	-- 0x1677
		when 005752 => D <= "11000011";	-- 0x1678
		when 005753 => D <= "01111110";	-- 0x1679
		when 005754 => D <= "00110110";	-- 0x167A
		when 005755 => D <= "11000011";	-- 0x167B
		when 005756 => D <= "01101110";	-- 0x167C
		when 005757 => D <= "00111111";	-- 0x167D
		when 005758 => D <= "11001001";	-- 0x167E
		when 005759 => D <= "11001101";	-- 0x167F
		when 005760 => D <= "00100010";	-- 0x1680
		when 005761 => D <= "00111100";	-- 0x1681
		when 005762 => D <= "11011010";	-- 0x1682
		when 005763 => D <= "01101110";	-- 0x1683
		when 005764 => D <= "00111111";	-- 0x1684
		when 005765 => D <= "01111100";	-- 0x1685
		when 005766 => D <= "10110101";	-- 0x1686
		when 005767 => D <= "11000010";	-- 0x1687
		when 005768 => D <= "10001110";	-- 0x1688
		when 005769 => D <= "00110110";	-- 0x1689
		when 005770 => D <= "10101111";	-- 0x168A
		when 005771 => D <= "11000011";	-- 0x168B
		when 005772 => D <= "10010000";	-- 0x168C
		when 005773 => D <= "00110110";	-- 0x168D
		when 005774 => D <= "00111110";	-- 0x168E
		when 005775 => D <= "11111111";	-- 0x168F
		when 005776 => D <= "00110010";	-- 0x1690
		when 005777 => D <= "00000011";	-- 0x1691
		when 005778 => D <= "10000000";	-- 0x1692
		when 005779 => D <= "11001001";	-- 0x1693
		when 005780 => D <= "00111010";	-- 0x1694
		when 005781 => D <= "00000011";	-- 0x1695
		when 005782 => D <= "10000000";	-- 0x1696
		when 005783 => D <= "10110111";	-- 0x1697
		when 005784 => D <= "11000010";	-- 0x1698
		when 005785 => D <= "10101010";	-- 0x1699
		when 005786 => D <= "00110110";	-- 0x169A
		when 005787 => D <= "11011101";	-- 0x169B
		when 005788 => D <= "01111110";	-- 0x169C
		when 005789 => D <= "00000000";	-- 0x169D
		when 005790 => D <= "10110111";	-- 0x169E
		when 005791 => D <= "11001010";	-- 0x169F
		when 005792 => D <= "10101010";	-- 0x16A0
		when 005793 => D <= "00110110";	-- 0x16A1
		when 005794 => D <= "11011101";	-- 0x16A2
		when 005795 => D <= "00100011";	-- 0x16A3
		when 005796 => D <= "11011101";	-- 0x16A4
		when 005797 => D <= "01111110";	-- 0x16A5
		when 005798 => D <= "00000000";	-- 0x16A6
		when 005799 => D <= "11000011";	-- 0x16A7
		when 005800 => D <= "10011110";	-- 0x16A8
		when 005801 => D <= "00110110";	-- 0x16A9
		when 005802 => D <= "11001001";	-- 0x16AA
		when 005803 => D <= "00111010";	-- 0x16AB
		when 005804 => D <= "00000011";	-- 0x16AC
		when 005805 => D <= "10000000";	-- 0x16AD
		when 005806 => D <= "10110111";	-- 0x16AE
		when 005807 => D <= "11001010";	-- 0x16AF
		when 005808 => D <= "11000001";	-- 0x16B0
		when 005809 => D <= "00110110";	-- 0x16B1
		when 005810 => D <= "11011101";	-- 0x16B2
		when 005811 => D <= "01111110";	-- 0x16B3
		when 005812 => D <= "00000000";	-- 0x16B4
		when 005813 => D <= "10110111";	-- 0x16B5
		when 005814 => D <= "11001010";	-- 0x16B6
		when 005815 => D <= "11000001";	-- 0x16B7
		when 005816 => D <= "00110110";	-- 0x16B8
		when 005817 => D <= "11011101";	-- 0x16B9
		when 005818 => D <= "00100011";	-- 0x16BA
		when 005819 => D <= "11011101";	-- 0x16BB
		when 005820 => D <= "01111110";	-- 0x16BC
		when 005821 => D <= "00000000";	-- 0x16BD
		when 005822 => D <= "11000011";	-- 0x16BE
		when 005823 => D <= "10110101";	-- 0x16BF
		when 005824 => D <= "00110110";	-- 0x16C0
		when 005825 => D <= "11001001";	-- 0x16C1
		when 005826 => D <= "11011101";	-- 0x16C2
		when 005827 => D <= "11100101";	-- 0x16C3
		when 005828 => D <= "11001101";	-- 0x16C4
		when 005829 => D <= "00100010";	-- 0x16C5
		when 005830 => D <= "00111100";	-- 0x16C6
		when 005831 => D <= "11011010";	-- 0x16C7
		when 005832 => D <= "01101110";	-- 0x16C8
		when 005833 => D <= "00111111";	-- 0x16C9
		when 005834 => D <= "01111101";	-- 0x16CA
		when 005835 => D <= "10110100";	-- 0x16CB
		when 005836 => D <= "11001010";	-- 0x16CC
		when 005837 => D <= "00000010";	-- 0x16CD
		when 005838 => D <= "00110111";	-- 0x16CE
		when 005839 => D <= "11001101";	-- 0x16CF
		when 005840 => D <= "11001100";	-- 0x16D0
		when 005841 => D <= "00100111";	-- 0x16D1
		when 005842 => D <= "11011101";	-- 0x16D2
		when 005843 => D <= "01111110";	-- 0x16D3
		when 005844 => D <= "00000000";	-- 0x16D4
		when 005845 => D <= "11111110";	-- 0x16D5
		when 005846 => D <= "01011011";	-- 0x16D6
		when 005847 => D <= "11000010";	-- 0x16D7
		when 005848 => D <= "11111011";	-- 0x16D8
		when 005849 => D <= "00110110";	-- 0x16D9
		when 005850 => D <= "11011101";	-- 0x16DA
		when 005851 => D <= "00100011";	-- 0x16DB
		when 005852 => D <= "11111110";	-- 0x16DC
		when 005853 => D <= "01011101";	-- 0x16DD
		when 005854 => D <= "11001010";	-- 0x16DE
		when 005855 => D <= "11110001";	-- 0x16DF
		when 005856 => D <= "00110110";	-- 0x16E0
		when 005857 => D <= "10110111";	-- 0x16E1
		when 005858 => D <= "11001010";	-- 0x16E2
		when 005859 => D <= "11110001";	-- 0x16E3
		when 005860 => D <= "00110110";	-- 0x16E4
		when 005861 => D <= "11001101";	-- 0x16E5
		when 005862 => D <= "00111011";	-- 0x16E6
		when 005863 => D <= "00111100";	-- 0x16E7
		when 005864 => D <= "11001101";	-- 0x16E8
		when 005865 => D <= "11001100";	-- 0x16E9
		when 005866 => D <= "00100111";	-- 0x16EA
		when 005867 => D <= "11011101";	-- 0x16EB
		when 005868 => D <= "01111110";	-- 0x16EC
		when 005869 => D <= "00000000";	-- 0x16ED
		when 005870 => D <= "11000011";	-- 0x16EE
		when 005871 => D <= "11011100";	-- 0x16EF
		when 005872 => D <= "00110110";	-- 0x16F0
		when 005873 => D <= "11111110";	-- 0x16F1
		when 005874 => D <= "01011101";	-- 0x16F2
		when 005875 => D <= "11000010";	-- 0x16F3
		when 005876 => D <= "11111000";	-- 0x16F4
		when 005877 => D <= "00110110";	-- 0x16F5
		when 005878 => D <= "11011101";	-- 0x16F6
		when 005879 => D <= "00100011";	-- 0x16F7
		when 005880 => D <= "11000011";	-- 0x16F8
		when 005881 => D <= "11111110";	-- 0x16F9
		when 005882 => D <= "00110110";	-- 0x16FA
		when 005883 => D <= "11000011";	-- 0x16FB
		when 005884 => D <= "01101110";	-- 0x16FC
		when 005885 => D <= "00111111";	-- 0x16FD
		when 005886 => D <= "11011101";	-- 0x16FE
		when 005887 => D <= "11100001";	-- 0x16FF
		when 005888 => D <= "00011000";	-- 0x1700
		when 005889 => D <= "11000000";	-- 0x1701
		when 005890 => D <= "11100001";	-- 0x1702
		when 005891 => D <= "11011010";	-- 0x1703
		when 005892 => D <= "01101110";	-- 0x1704
		when 005893 => D <= "00111111";	-- 0x1705
		when 005894 => D <= "11001101";	-- 0x1706
		when 005895 => D <= "11001100";	-- 0x1707
		when 005896 => D <= "00100111";	-- 0x1708
		when 005897 => D <= "11001101";	-- 0x1709
		when 005898 => D <= "10110100";	-- 0x170A
		when 005899 => D <= "00110111";	-- 0x170B
		when 005900 => D <= "11001001";	-- 0x170C
		when 005901 => D <= "00111110";	-- 0x170D
		when 005902 => D <= "00000001";	-- 0x170E
		when 005903 => D <= "00110010";	-- 0x170F
		when 005904 => D <= "00000100";	-- 0x1710
		when 005905 => D <= "10000000";	-- 0x1711
		when 005906 => D <= "11001001";	-- 0x1712
		when 005907 => D <= "10101111";	-- 0x1713
		when 005908 => D <= "00011000";	-- 0x1714
		when 005909 => D <= "11111001";	-- 0x1715
		when 005910 => D <= "00111010";	-- 0x1716
		when 005911 => D <= "00000010";	-- 0x1717
		when 005912 => D <= "10000000";	-- 0x1718
		when 005913 => D <= "10110111";	-- 0x1719
		when 005914 => D <= "11001010";	-- 0x171A
		when 005915 => D <= "00100000";	-- 0x171B
		when 005916 => D <= "00110111";	-- 0x171C
		when 005917 => D <= "11000011";	-- 0x171D
		when 005918 => D <= "01101110";	-- 0x171E
		when 005919 => D <= "00111111";	-- 0x171F
		when 005920 => D <= "11001101";	-- 0x1720
		when 005921 => D <= "11001100";	-- 0x1721
		when 005922 => D <= "00100111";	-- 0x1722
		when 005923 => D <= "11011101";	-- 0x1723
		when 005924 => D <= "01111110";	-- 0x1724
		when 005925 => D <= "00000000";	-- 0x1725
		when 005926 => D <= "10110111";	-- 0x1726
		when 005927 => D <= "11000010";	-- 0x1727
		when 005928 => D <= "01000101";	-- 0x1728
		when 005929 => D <= "00110111";	-- 0x1729
		when 005930 => D <= "00100001";	-- 0x172A
		when 005931 => D <= "01101001";	-- 0x172B
		when 005932 => D <= "00110111";	-- 0x172C
		when 005933 => D <= "11001101";	-- 0x172D
		when 005934 => D <= "10110010";	-- 0x172E
		when 005935 => D <= "00111110";	-- 0x172F
		when 005936 => D <= "11001101";	-- 0x1730
		when 005937 => D <= "00101001";	-- 0x1731
		when 005938 => D <= "00100000";	-- 0x1732
		when 005939 => D <= "01001111";	-- 0x1733
		when 005940 => D <= "11001101";	-- 0x1734
		when 005941 => D <= "10110111";	-- 0x1735
		when 005942 => D <= "00110000";	-- 0x1736
		when 005943 => D <= "11111110";	-- 0x1737
		when 005944 => D <= "01001010";	-- 0x1738
		when 005945 => D <= "11000010";	-- 0x1739
		when 005946 => D <= "00111111";	-- 0x173A
		when 005947 => D <= "00110111";	-- 0x173B
		when 005948 => D <= "11001101";	-- 0x173C
		when 005949 => D <= "00000111";	-- 0x173D
		when 005950 => D <= "00111110";	-- 0x173E
		when 005951 => D <= "11001101";	-- 0x173F
		when 005952 => D <= "11101111";	-- 0x1740
		when 005953 => D <= "00110000";	-- 0x1741
		when 005954 => D <= "11000011";	-- 0x1742
		when 005955 => D <= "01101000";	-- 0x1743
		when 005956 => D <= "00110111";	-- 0x1744
		when 005957 => D <= "11111101";	-- 0x1745
		when 005958 => D <= "00100001";	-- 0x1746
		when 005959 => D <= "01001111";	-- 0x1747
		when 005960 => D <= "10000011";	-- 0x1748
		when 005961 => D <= "11011101";	-- 0x1749
		when 005962 => D <= "11100101";	-- 0x174A
		when 005963 => D <= "11001101";	-- 0x174B
		when 005964 => D <= "00110101";	-- 0x174C
		when 005965 => D <= "00101010";	-- 0x174D
		when 005966 => D <= "11011101";	-- 0x174E
		when 005967 => D <= "11100001";	-- 0x174F
		when 005968 => D <= "11011010";	-- 0x1750
		when 005969 => D <= "01101000";	-- 0x1751
		when 005970 => D <= "00110111";	-- 0x1752
		when 005971 => D <= "11111110";	-- 0x1753
		when 005972 => D <= "00000010";	-- 0x1754
		when 005973 => D <= "11000010";	-- 0x1755
		when 005974 => D <= "01100101";	-- 0x1756
		when 005975 => D <= "00110111";	-- 0x1757
		when 005976 => D <= "11011101";	-- 0x1758
		when 005977 => D <= "11100101";	-- 0x1759
		when 005978 => D <= "11001101";	-- 0x175A
		when 005979 => D <= "00100011";	-- 0x175B
		when 005980 => D <= "00110100";	-- 0x175C
		when 005981 => D <= "11011101";	-- 0x175D
		when 005982 => D <= "11100001";	-- 0x175E
		when 005983 => D <= "11001101";	-- 0x175F
		when 005984 => D <= "11100011";	-- 0x1760
		when 005985 => D <= "00101010";	-- 0x1761
		when 005986 => D <= "11000011";	-- 0x1762
		when 005987 => D <= "01101000";	-- 0x1763
		when 005988 => D <= "00110111";	-- 0x1764
		when 005989 => D <= "11001101";	-- 0x1765
		when 005990 => D <= "11100011";	-- 0x1766
		when 005991 => D <= "00101010";	-- 0x1767
		when 005992 => D <= "11001001";	-- 0x1768
		when 005993 => D <= "01000001";	-- 0x1769
		when 005994 => D <= "01101100";	-- 0x176A
		when 005995 => D <= "01101100";	-- 0x176B
		when 005996 => D <= "01100101";	-- 0x176C
		when 005997 => D <= "01110011";	-- 0x176D
		when 005998 => D <= "00100000";	-- 0x176E
		when 005999 => D <= "00111111";	-- 0x176F
		when 006000 => D <= "00100000";	-- 0x1770
		when 006001 => D <= "01001010";	-- 0x1771
		when 006002 => D <= "00111101";	-- 0x1772
		when 006003 => D <= "01001010";	-- 0x1773
		when 006004 => D <= "01000001";	-- 0x1774
		when 006005 => D <= "00100000";	-- 0x1775
		when 006006 => D <= "00000000";	-- 0x1776
		when 006007 => D <= "11001101";	-- 0x1777
		when 006008 => D <= "00100010";	-- 0x1778
		when 006009 => D <= "00111100";	-- 0x1779
		when 006010 => D <= "11011010";	-- 0x177A
		when 006011 => D <= "01101110";	-- 0x177B
		when 006012 => D <= "00111111";	-- 0x177C
		when 006013 => D <= "01111100";	-- 0x177D
		when 006014 => D <= "10110101";	-- 0x177E
		when 006015 => D <= "00101000";	-- 0x177F
		when 006016 => D <= "00101100";	-- 0x1780
		when 006017 => D <= "00101011";	-- 0x1781
		when 006018 => D <= "11100101";	-- 0x1782
		when 006019 => D <= "11011101";	-- 0x1783
		when 006020 => D <= "11100101";	-- 0x1784
		when 006021 => D <= "11001101";	-- 0x1785
		when 006022 => D <= "11001100";	-- 0x1786
		when 006023 => D <= "00100111";	-- 0x1787
		when 006024 => D <= "11111110";	-- 0x1788
		when 006025 => D <= "01011011";	-- 0x1789
		when 006026 => D <= "11000010";	-- 0x178A
		when 006027 => D <= "10101000";	-- 0x178B
		when 006028 => D <= "00110111";	-- 0x178C
		when 006029 => D <= "11011101";	-- 0x178D
		when 006030 => D <= "00100011";	-- 0x178E
		when 006031 => D <= "11001101";	-- 0x178F
		when 006032 => D <= "00111011";	-- 0x1790
		when 006033 => D <= "00111100";	-- 0x1791
		when 006034 => D <= "11001101";	-- 0x1792
		when 006035 => D <= "11001100";	-- 0x1793
		when 006036 => D <= "00100111";	-- 0x1794
		when 006037 => D <= "11011101";	-- 0x1795
		when 006038 => D <= "01111110";	-- 0x1796
		when 006039 => D <= "00000000";	-- 0x1797
		when 006040 => D <= "11111110";	-- 0x1798
		when 006041 => D <= "01011101";	-- 0x1799
		when 006042 => D <= "11001010";	-- 0x179A
		when 006043 => D <= "10100001";	-- 0x179B
		when 006044 => D <= "00110111";	-- 0x179C
		when 006045 => D <= "10110111";	-- 0x179D
		when 006046 => D <= "11000010";	-- 0x179E
		when 006047 => D <= "10001111";	-- 0x179F
		when 006048 => D <= "00110111";	-- 0x17A0
		when 006049 => D <= "11111110";	-- 0x17A1
		when 006050 => D <= "01011101";	-- 0x17A2
		when 006051 => D <= "11000010";	-- 0x17A3
		when 006052 => D <= "10101000";	-- 0x17A4
		when 006053 => D <= "00110111";	-- 0x17A5
		when 006054 => D <= "11011101";	-- 0x17A6
		when 006055 => D <= "00100011";	-- 0x17A7
		when 006056 => D <= "11011101";	-- 0x17A8
		when 006057 => D <= "11100001";	-- 0x17A9
		when 006058 => D <= "11100001";	-- 0x17AA
		when 006059 => D <= "00011000";	-- 0x17AB
		when 006060 => D <= "11010000";	-- 0x17AC
		when 006061 => D <= "11001101";	-- 0x17AD
		when 006062 => D <= "11001100";	-- 0x17AE
		when 006063 => D <= "00100111";	-- 0x17AF
		when 006064 => D <= "11001101";	-- 0x17B0
		when 006065 => D <= "10110100";	-- 0x17B1
		when 006066 => D <= "00110111";	-- 0x17B2
		when 006067 => D <= "11001001";	-- 0x17B3
		when 006068 => D <= "11011101";	-- 0x17B4
		when 006069 => D <= "01111110";	-- 0x17B5
		when 006070 => D <= "00000000";	-- 0x17B6
		when 006071 => D <= "11111110";	-- 0x17B7
		when 006072 => D <= "01011011";	-- 0x17B8
		when 006073 => D <= "11000000";	-- 0x17B9
		when 006074 => D <= "11011101";	-- 0x17BA
		when 006075 => D <= "00100011";	-- 0x17BB
		when 006076 => D <= "11011101";	-- 0x17BC
		when 006077 => D <= "01111110";	-- 0x17BD
		when 006078 => D <= "00000000";	-- 0x17BE
		when 006079 => D <= "11111110";	-- 0x17BF
		when 006080 => D <= "01011011";	-- 0x17C0
		when 006081 => D <= "11000010";	-- 0x17C1
		when 006082 => D <= "11000111";	-- 0x17C2
		when 006083 => D <= "00110111";	-- 0x17C3
		when 006084 => D <= "11001101";	-- 0x17C4
		when 006085 => D <= "10110100";	-- 0x17C5
		when 006086 => D <= "00110111";	-- 0x17C6
		when 006087 => D <= "11011101";	-- 0x17C7
		when 006088 => D <= "01111110";	-- 0x17C8
		when 006089 => D <= "00000000";	-- 0x17C9
		when 006090 => D <= "11011101";	-- 0x17CA
		when 006091 => D <= "00100011";	-- 0x17CB
		when 006092 => D <= "11111110";	-- 0x17CC
		when 006093 => D <= "01011101";	-- 0x17CD
		when 006094 => D <= "11001010";	-- 0x17CE
		when 006095 => D <= "11010101";	-- 0x17CF
		when 006096 => D <= "00110111";	-- 0x17D0
		when 006097 => D <= "10110111";	-- 0x17D1
		when 006098 => D <= "11000010";	-- 0x17D2
		when 006099 => D <= "10111100";	-- 0x17D3
		when 006100 => D <= "00110111";	-- 0x17D4
		when 006101 => D <= "10110111";	-- 0x17D5
		when 006102 => D <= "11000010";	-- 0x17D6
		when 006103 => D <= "11011011";	-- 0x17D7
		when 006104 => D <= "00110111";	-- 0x17D8
		when 006105 => D <= "11011101";	-- 0x17D9
		when 006106 => D <= "00101011";	-- 0x17DA
		when 006107 => D <= "11001001";	-- 0x17DB
		when 006108 => D <= "00111010";	-- 0x17DC
		when 006109 => D <= "00000010";	-- 0x17DD
		when 006110 => D <= "10000000";	-- 0x17DE
		when 006111 => D <= "11111110";	-- 0x17DF
		when 006112 => D <= "11111111";	-- 0x17E0
		when 006113 => D <= "11000010";	-- 0x17E1
		when 006114 => D <= "11101011";	-- 0x17E2
		when 006115 => D <= "00110111";	-- 0x17E3
		when 006116 => D <= "10101111";	-- 0x17E4
		when 006117 => D <= "00110010";	-- 0x17E5
		when 006118 => D <= "00000010";	-- 0x17E6
		when 006119 => D <= "10000000";	-- 0x17E7
		when 006120 => D <= "11000011";	-- 0x17E8
		when 006121 => D <= "11101110";	-- 0x17E9
		when 006122 => D <= "00110111";	-- 0x17EA
		when 006123 => D <= "11000011";	-- 0x17EB
		when 006124 => D <= "01101110";	-- 0x17EC
		when 006125 => D <= "00111111";	-- 0x17ED
		when 006126 => D <= "11001001";	-- 0x17EE
		when 006127 => D <= "11001101";	-- 0x17EF
		when 006128 => D <= "11001100";	-- 0x17F0
		when 006129 => D <= "00100111";	-- 0x17F1
		when 006130 => D <= "11011101";	-- 0x17F2
		when 006131 => D <= "01111110";	-- 0x17F3
		when 006132 => D <= "00000000";	-- 0x17F4
		when 006133 => D <= "11111110";	-- 0x17F5
		when 006134 => D <= "00100010";	-- 0x17F6
		when 006135 => D <= "11000010";	-- 0x17F7
		when 006136 => D <= "00010110";	-- 0x17F8
		when 006137 => D <= "00111000";	-- 0x17F9
		when 006138 => D <= "11011101";	-- 0x17FA
		when 006139 => D <= "00100011";	-- 0x17FB
		when 006140 => D <= "11111110";	-- 0x17FC
		when 006141 => D <= "00100000";	-- 0x17FD
		when 006142 => D <= "11001010";	-- 0x17FE
		when 006143 => D <= "00010011";	-- 0x17FF
		when 006144 => D <= "00111000";	-- 0x1800
		when 006145 => D <= "10110111";	-- 0x1801
		when 006146 => D <= "11001010";	-- 0x1802
		when 006147 => D <= "00010011";	-- 0x1803
		when 006148 => D <= "00111000";	-- 0x1804
		when 006149 => D <= "11011101";	-- 0x1805
		when 006150 => D <= "01001110";	-- 0x1806
		when 006151 => D <= "00000000";	-- 0x1807
		when 006152 => D <= "11001101";	-- 0x1808
		when 006153 => D <= "10110111";	-- 0x1809
		when 006154 => D <= "00110000";	-- 0x180A
		when 006155 => D <= "11011101";	-- 0x180B
		when 006156 => D <= "00100011";	-- 0x180C
		when 006157 => D <= "11011101";	-- 0x180D
		when 006158 => D <= "01111110";	-- 0x180E
		when 006159 => D <= "00000000";	-- 0x180F
		when 006160 => D <= "11000011";	-- 0x1810
		when 006161 => D <= "11111100";	-- 0x1811
		when 006162 => D <= "00110111";	-- 0x1812
		when 006163 => D <= "11000011";	-- 0x1813
		when 006164 => D <= "01011100";	-- 0x1814
		when 006165 => D <= "00111000";	-- 0x1815
		when 006166 => D <= "11111110";	-- 0x1816
		when 006167 => D <= "01011011";	-- 0x1817
		when 006168 => D <= "11000010";	-- 0x1818
		when 006169 => D <= "01010110";	-- 0x1819
		when 006170 => D <= "00111000";	-- 0x181A
		when 006171 => D <= "11011101";	-- 0x181B
		when 006172 => D <= "00100011";	-- 0x181C
		when 006173 => D <= "11011101";	-- 0x181D
		when 006174 => D <= "01111110";	-- 0x181E
		when 006175 => D <= "00000000";	-- 0x181F
		when 006176 => D <= "11111110";	-- 0x1820
		when 006177 => D <= "01011101";	-- 0x1821
		when 006178 => D <= "11001010";	-- 0x1822
		when 006179 => D <= "01001100";	-- 0x1823
		when 006180 => D <= "00111000";	-- 0x1824
		when 006181 => D <= "10110111";	-- 0x1825
		when 006182 => D <= "11001010";	-- 0x1826
		when 006183 => D <= "01001100";	-- 0x1827
		when 006184 => D <= "00111000";	-- 0x1828
		when 006185 => D <= "11111110";	-- 0x1829
		when 006186 => D <= "01011011";	-- 0x182A
		when 006187 => D <= "11000010";	-- 0x182B
		when 006188 => D <= "00111110";	-- 0x182C
		when 006189 => D <= "00111000";	-- 0x182D
		when 006190 => D <= "00001110";	-- 0x182E
		when 006191 => D <= "01011011";	-- 0x182F
		when 006192 => D <= "11001101";	-- 0x1830
		when 006193 => D <= "10110111";	-- 0x1831
		when 006194 => D <= "00110000";	-- 0x1832
		when 006195 => D <= "11001101";	-- 0x1833
		when 006196 => D <= "11101111";	-- 0x1834
		when 006197 => D <= "00110111";	-- 0x1835
		when 006198 => D <= "00001110";	-- 0x1836
		when 006199 => D <= "01011101";	-- 0x1837
		when 006200 => D <= "11001101";	-- 0x1838
		when 006201 => D <= "10110111";	-- 0x1839
		when 006202 => D <= "00110000";	-- 0x183A
		when 006203 => D <= "11000011";	-- 0x183B
		when 006204 => D <= "01000110";	-- 0x183C
		when 006205 => D <= "00111000";	-- 0x183D
		when 006206 => D <= "11011101";	-- 0x183E
		when 006207 => D <= "01001110";	-- 0x183F
		when 006208 => D <= "00000000";	-- 0x1840
		when 006209 => D <= "11001101";	-- 0x1841
		when 006210 => D <= "10110111";	-- 0x1842
		when 006211 => D <= "00110000";	-- 0x1843
		when 006212 => D <= "11011101";	-- 0x1844
		when 006213 => D <= "00100011";	-- 0x1845
		when 006214 => D <= "11011101";	-- 0x1846
		when 006215 => D <= "01111110";	-- 0x1847
		when 006216 => D <= "00000000";	-- 0x1848
		when 006217 => D <= "11000011";	-- 0x1849
		when 006218 => D <= "00100000";	-- 0x184A
		when 006219 => D <= "00111000";	-- 0x184B
		when 006220 => D <= "11111110";	-- 0x184C
		when 006221 => D <= "01011101";	-- 0x184D
		when 006222 => D <= "11000010";	-- 0x184E
		when 006223 => D <= "01010011";	-- 0x184F
		when 006224 => D <= "00111000";	-- 0x1850
		when 006225 => D <= "11011101";	-- 0x1851
		when 006226 => D <= "00100011";	-- 0x1852
		when 006227 => D <= "11000011";	-- 0x1853
		when 006228 => D <= "01011100";	-- 0x1854
		when 006229 => D <= "00111000";	-- 0x1855
		when 006230 => D <= "11001101";	-- 0x1856
		when 006231 => D <= "00100010";	-- 0x1857
		when 006232 => D <= "00111100";	-- 0x1858
		when 006233 => D <= "11001101";	-- 0x1859
		when 006234 => D <= "00001111";	-- 0x185A
		when 006235 => D <= "00101010";	-- 0x185B
		when 006236 => D <= "11001001";	-- 0x185C
		when 006237 => D <= "11001101";	-- 0x185D
		when 006238 => D <= "11101111";	-- 0x185E
		when 006239 => D <= "00110111";	-- 0x185F
		when 006240 => D <= "11001101";	-- 0x1860
		when 006241 => D <= "11101111";	-- 0x1861
		when 006242 => D <= "00110000";	-- 0x1862
		when 006243 => D <= "11001001";	-- 0x1863
		when 006244 => D <= "11001101";	-- 0x1864
		when 006245 => D <= "00100010";	-- 0x1865
		when 006246 => D <= "00111100";	-- 0x1866
		when 006247 => D <= "11011010";	-- 0x1867
		when 006248 => D <= "01101110";	-- 0x1868
		when 006249 => D <= "00111111";	-- 0x1869
		when 006250 => D <= "01001101";	-- 0x186A
		when 006251 => D <= "11001101";	-- 0x186B
		when 006252 => D <= "10110111";	-- 0x186C
		when 006253 => D <= "00110000";	-- 0x186D
		when 006254 => D <= "11001001";	-- 0x186E
		when 006255 => D <= "11001101";	-- 0x186F
		when 006256 => D <= "00100010";	-- 0x1870
		when 006257 => D <= "00111100";	-- 0x1871
		when 006258 => D <= "11011010";	-- 0x1872
		when 006259 => D <= "01101110";	-- 0x1873
		when 006260 => D <= "00111111";	-- 0x1874
		when 006261 => D <= "11100101";	-- 0x1875
		when 006262 => D <= "11001101";	-- 0x1876
		when 006263 => D <= "00100010";	-- 0x1877
		when 006264 => D <= "00111100";	-- 0x1878
		when 006265 => D <= "11011010";	-- 0x1879
		when 006266 => D <= "01101110";	-- 0x187A
		when 006267 => D <= "00111111";	-- 0x187B
		when 006268 => D <= "11010001";	-- 0x187C
		when 006269 => D <= "01001011";	-- 0x187D
		when 006270 => D <= "11101101";	-- 0x187E
		when 006271 => D <= "01101001";	-- 0x187F
		when 006272 => D <= "11001001";	-- 0x1880
		when 006273 => D <= "11001001";	-- 0x1881
		when 006274 => D <= "11001101";	-- 0x1882
		when 006275 => D <= "00111010";	-- 0x1883
		when 006276 => D <= "00100100";	-- 0x1884
		when 006277 => D <= "00100001";	-- 0x1885
		when 006278 => D <= "01011010";	-- 0x1886
		when 006279 => D <= "00000000";	-- 0x1887
		when 006280 => D <= "00100010";	-- 0x1888
		when 006281 => D <= "00111011";	-- 0x1889
		when 006282 => D <= "10000000";	-- 0x188A
		when 006283 => D <= "00100001";	-- 0x188B
		when 006284 => D <= "00000000";	-- 0x188C
		when 006285 => D <= "00000001";	-- 0x188D
		when 006286 => D <= "11001101";	-- 0x188E
		when 006287 => D <= "00010100";	-- 0x188F
		when 006288 => D <= "00100101";	-- 0x1890
		when 006289 => D <= "11101011";	-- 0x1891
		when 006290 => D <= "00100001";	-- 0x1892
		when 006291 => D <= "00000000";	-- 0x1893
		when 006292 => D <= "00000001";	-- 0x1894
		when 006293 => D <= "11001101";	-- 0x1895
		when 006294 => D <= "00010100";	-- 0x1896
		when 006295 => D <= "00100101";	-- 0x1897
		when 006296 => D <= "11000011";	-- 0x1898
		when 006297 => D <= "11010111";	-- 0x1899
		when 006298 => D <= "00111000";	-- 0x189A
		when 006299 => D <= "11001101";	-- 0x189B
		when 006300 => D <= "00111010";	-- 0x189C
		when 006301 => D <= "00100100";	-- 0x189D
		when 006302 => D <= "11001101";	-- 0x189E
		when 006303 => D <= "00100010";	-- 0x189F
		when 006304 => D <= "00111100";	-- 0x18A0
		when 006305 => D <= "11011010";	-- 0x18A1
		when 006306 => D <= "01101110";	-- 0x18A2
		when 006307 => D <= "00111111";	-- 0x18A3
		when 006308 => D <= "11001101";	-- 0x18A4
		when 006309 => D <= "00010100";	-- 0x18A5
		when 006310 => D <= "00100101";	-- 0x18A6
		when 006311 => D <= "11101101";	-- 0x18A7
		when 006312 => D <= "01011011";	-- 0x18A8
		when 006313 => D <= "00111001";	-- 0x18A9
		when 006314 => D <= "10000000";	-- 0x18AA
		when 006315 => D <= "00011000";	-- 0x18AB
		when 006316 => D <= "00101010";	-- 0x18AC
		when 006317 => D <= "11001101";	-- 0x18AD
		when 006318 => D <= "00111010";	-- 0x18AE
		when 006319 => D <= "00100100";	-- 0x18AF
		when 006320 => D <= "11001101";	-- 0x18B0
		when 006321 => D <= "00100010";	-- 0x18B1
		when 006322 => D <= "00111100";	-- 0x18B2
		when 006323 => D <= "11011010";	-- 0x18B3
		when 006324 => D <= "01101110";	-- 0x18B4
		when 006325 => D <= "00111111";	-- 0x18B5
		when 006326 => D <= "11001101";	-- 0x18B6
		when 006327 => D <= "00010100";	-- 0x18B7
		when 006328 => D <= "00100101";	-- 0x18B8
		when 006329 => D <= "11101011";	-- 0x18B9
		when 006330 => D <= "00101010";	-- 0x18BA
		when 006331 => D <= "00110111";	-- 0x18BB
		when 006332 => D <= "10000000";	-- 0x18BC
		when 006333 => D <= "00011000";	-- 0x18BD
		when 006334 => D <= "00011000";	-- 0x18BE
		when 006335 => D <= "11001101";	-- 0x18BF
		when 006336 => D <= "00111010";	-- 0x18C0
		when 006337 => D <= "00100100";	-- 0x18C1
		when 006338 => D <= "11001101";	-- 0x18C2
		when 006339 => D <= "00100010";	-- 0x18C3
		when 006340 => D <= "00111100";	-- 0x18C4
		when 006341 => D <= "11011010";	-- 0x18C5
		when 006342 => D <= "01101110";	-- 0x18C6
		when 006343 => D <= "00111111";	-- 0x18C7
		when 006344 => D <= "11001101";	-- 0x18C8
		when 006345 => D <= "00010100";	-- 0x18C9
		when 006346 => D <= "00100101";	-- 0x18CA
		when 006347 => D <= "11100101";	-- 0x18CB
		when 006348 => D <= "11001101";	-- 0x18CC
		when 006349 => D <= "00100010";	-- 0x18CD
		when 006350 => D <= "00111100";	-- 0x18CE
		when 006351 => D <= "11011010";	-- 0x18CF
		when 006352 => D <= "01101110";	-- 0x18D0
		when 006353 => D <= "00111111";	-- 0x18D1
		when 006354 => D <= "11001101";	-- 0x18D2
		when 006355 => D <= "00010100";	-- 0x18D3
		when 006356 => D <= "00100101";	-- 0x18D4
		when 006357 => D <= "11010001";	-- 0x18D5
		when 006358 => D <= "11101011";	-- 0x18D6
		when 006359 => D <= "00100010";	-- 0x18D7
		when 006360 => D <= "00110111";	-- 0x18D8
		when 006361 => D <= "10000000";	-- 0x18D9
		when 006362 => D <= "11101101";	-- 0x18DA
		when 006363 => D <= "01010011";	-- 0x18DB
		when 006364 => D <= "00111001";	-- 0x18DC
		when 006365 => D <= "10000000";	-- 0x18DD
		when 006366 => D <= "11000011";	-- 0x18DE
		when 006367 => D <= "10010011";	-- 0x18DF
		when 006368 => D <= "00100100";	-- 0x18E0
		when 006369 => D <= "11001101";	-- 0x18E1
		when 006370 => D <= "00100010";	-- 0x18E2
		when 006371 => D <= "00111100";	-- 0x18E3
		when 006372 => D <= "11011010";	-- 0x18E4
		when 006373 => D <= "01101110";	-- 0x18E5
		when 006374 => D <= "00111111";	-- 0x18E6
		when 006375 => D <= "11000011";	-- 0x18E7
		when 006376 => D <= "00011000";	-- 0x18E8
		when 006377 => D <= "00100100";	-- 0x18E9
		when 006378 => D <= "11001101";	-- 0x18EA
		when 006379 => D <= "00010001";	-- 0x18EB
		when 006380 => D <= "00100001";	-- 0x18EC
		when 006381 => D <= "11001001";	-- 0x18ED
		when 006382 => D <= "11001101";	-- 0x18EE
		when 006383 => D <= "00100010";	-- 0x18EF
		when 006384 => D <= "00111100";	-- 0x18F0
		when 006385 => D <= "11011010";	-- 0x18F1
		when 006386 => D <= "01101110";	-- 0x18F2
		when 006387 => D <= "00111111";	-- 0x18F3
		when 006388 => D <= "01111101";	-- 0x18F4
		when 006389 => D <= "10110111";	-- 0x18F5
		when 006390 => D <= "11000010";	-- 0x18F6
		when 006391 => D <= "00000011";	-- 0x18F7
		when 006392 => D <= "00111001";	-- 0x18F8
		when 006393 => D <= "11001101";	-- 0x18F9
		when 006394 => D <= "01000010";	-- 0x18FA
		when 006395 => D <= "00100010";	-- 0x18FB
		when 006396 => D <= "10101111";	-- 0x18FC
		when 006397 => D <= "00110010";	-- 0x18FD
		when 006398 => D <= "00101001";	-- 0x18FE
		when 006399 => D <= "10000000";	-- 0x18FF
		when 006400 => D <= "11000011";	-- 0x1900
		when 006401 => D <= "00010001";	-- 0x1901
		when 006402 => D <= "00111001";	-- 0x1902
		when 006403 => D <= "01111101";	-- 0x1903
		when 006404 => D <= "11111110";	-- 0x1904
		when 006405 => D <= "00000001";	-- 0x1905
		when 006406 => D <= "11000010";	-- 0x1906
		when 006407 => D <= "00010001";	-- 0x1907
		when 006408 => D <= "00111001";	-- 0x1908
		when 006409 => D <= "11001101";	-- 0x1909
		when 006410 => D <= "01000110";	-- 0x190A
		when 006411 => D <= "00100010";	-- 0x190B
		when 006412 => D <= "00111110";	-- 0x190C
		when 006413 => D <= "00000001";	-- 0x190D
		when 006414 => D <= "00110010";	-- 0x190E
		when 006415 => D <= "00101001";	-- 0x190F
		when 006416 => D <= "10000000";	-- 0x1910
		when 006417 => D <= "11001001";	-- 0x1911
		when 006418 => D <= "00111110";	-- 0x1912
		when 006419 => D <= "00000001";	-- 0x1913
		when 006420 => D <= "00110010";	-- 0x1914
		when 006421 => D <= "00110110";	-- 0x1915
		when 006422 => D <= "10000000";	-- 0x1916
		when 006423 => D <= "11001101";	-- 0x1917
		when 006424 => D <= "00010001";	-- 0x1918
		when 006425 => D <= "00100001";	-- 0x1919
		when 006426 => D <= "11001001";	-- 0x191A
		when 006427 => D <= "11001101";	-- 0x191B
		when 006428 => D <= "00010001";	-- 0x191C
		when 006429 => D <= "00100001";	-- 0x191D
		when 006430 => D <= "11001101";	-- 0x191E
		when 006431 => D <= "11111101";	-- 0x191F
		when 006432 => D <= "00100011";	-- 0x1920
		when 006433 => D <= "11001001";	-- 0x1921
		when 006434 => D <= "11001101";	-- 0x1922
		when 006435 => D <= "00100010";	-- 0x1923
		when 006436 => D <= "00111100";	-- 0x1924
		when 006437 => D <= "11011010";	-- 0x1925
		when 006438 => D <= "01101110";	-- 0x1926
		when 006439 => D <= "00111111";	-- 0x1927
		when 006440 => D <= "01111101";	-- 0x1928
		when 006441 => D <= "00110010";	-- 0x1929
		when 006442 => D <= "00100111";	-- 0x192A
		when 006443 => D <= "10000000";	-- 0x192B
		when 006444 => D <= "00110010";	-- 0x192C
		when 006445 => D <= "00101000";	-- 0x192D
		when 006446 => D <= "10000000";	-- 0x192E
		when 006447 => D <= "11001101";	-- 0x192F
		when 006448 => D <= "00100010";	-- 0x1930
		when 006449 => D <= "00111100";	-- 0x1931
		when 006450 => D <= "11011010";	-- 0x1932
		when 006451 => D <= "01101110";	-- 0x1933
		when 006452 => D <= "00111111";	-- 0x1934
		when 006453 => D <= "01111101";	-- 0x1935
		when 006454 => D <= "00110010";	-- 0x1936
		when 006455 => D <= "00100101";	-- 0x1937
		when 006456 => D <= "10000000";	-- 0x1938
		when 006457 => D <= "00110010";	-- 0x1939
		when 006458 => D <= "00100110";	-- 0x193A
		when 006459 => D <= "10000000";	-- 0x193B
		when 006460 => D <= "11001001";	-- 0x193C
		when 006461 => D <= "11001101";	-- 0x193D
		when 006462 => D <= "00100010";	-- 0x193E
		when 006463 => D <= "00111100";	-- 0x193F
		when 006464 => D <= "11011010";	-- 0x1940
		when 006465 => D <= "01101110";	-- 0x1941
		when 006466 => D <= "00111111";	-- 0x1942
		when 006467 => D <= "11100101";	-- 0x1943
		when 006468 => D <= "11001101";	-- 0x1944
		when 006469 => D <= "00100010";	-- 0x1945
		when 006470 => D <= "00111100";	-- 0x1946
		when 006471 => D <= "11011010";	-- 0x1947
		when 006472 => D <= "01101110";	-- 0x1948
		when 006473 => D <= "00111111";	-- 0x1949
		when 006474 => D <= "11010001";	-- 0x194A
		when 006475 => D <= "01111101";	-- 0x194B
		when 006476 => D <= "00010010";	-- 0x194C
		when 006477 => D <= "11001001";	-- 0x194D
		when 006478 => D <= "11001101";	-- 0x194E
		when 006479 => D <= "11001100";	-- 0x194F
		when 006480 => D <= "00100111";	-- 0x1950
		when 006481 => D <= "11111101";	-- 0x1951
		when 006482 => D <= "00100001";	-- 0x1952
		when 006483 => D <= "01001111";	-- 0x1953
		when 006484 => D <= "10000011";	-- 0x1954
		when 006485 => D <= "11001101";	-- 0x1955
		when 006486 => D <= "00110101";	-- 0x1956
		when 006487 => D <= "00101010";	-- 0x1957
		when 006488 => D <= "11011010";	-- 0x1958
		when 006489 => D <= "10101011";	-- 0x1959
		when 006490 => D <= "00111001";	-- 0x195A
		when 006491 => D <= "11011101";	-- 0x195B
		when 006492 => D <= "11100101";	-- 0x195C
		when 006493 => D <= "11111110";	-- 0x195D
		when 006494 => D <= "00000001";	-- 0x195E
		when 006495 => D <= "11000010";	-- 0x195F
		when 006496 => D <= "01101011";	-- 0x1960
		when 006497 => D <= "00111001";	-- 0x1961
		when 006498 => D <= "11001101";	-- 0x1962
		when 006499 => D <= "00001111";	-- 0x1963
		when 006500 => D <= "00101010";	-- 0x1964
		when 006501 => D <= "11001101";	-- 0x1965
		when 006502 => D <= "11101111";	-- 0x1966
		when 006503 => D <= "00110000";	-- 0x1967
		when 006504 => D <= "11000011";	-- 0x1968
		when 006505 => D <= "10100110";	-- 0x1969
		when 006506 => D <= "00111001";	-- 0x196A
		when 006507 => D <= "11111110";	-- 0x196B
		when 006508 => D <= "00000010";	-- 0x196C
		when 006509 => D <= "11000010";	-- 0x196D
		when 006510 => D <= "10100110";	-- 0x196E
		when 006511 => D <= "00111001";	-- 0x196F
		when 006512 => D <= "11100101";	-- 0x1970
		when 006513 => D <= "11011101";	-- 0x1971
		when 006514 => D <= "11100001";	-- 0x1972
		when 006515 => D <= "11011101";	-- 0x1973
		when 006516 => D <= "11100101";	-- 0x1974
		when 006517 => D <= "11111101";	-- 0x1975
		when 006518 => D <= "00100001";	-- 0x1976
		when 006519 => D <= "10000111";	-- 0x1977
		when 006520 => D <= "00110001";	-- 0x1978
		when 006521 => D <= "11001101";	-- 0x1979
		when 006522 => D <= "11001100";	-- 0x197A
		when 006523 => D <= "00100111";	-- 0x197B
		when 006524 => D <= "11001101";	-- 0x197C
		when 006525 => D <= "00110101";	-- 0x197D
		when 006526 => D <= "00101010";	-- 0x197E
		when 006527 => D <= "11010010";	-- 0x197F
		when 006528 => D <= "10000100";	-- 0x1980
		when 006529 => D <= "00111001";	-- 0x1981
		when 006530 => D <= "00101110";	-- 0x1982
		when 006531 => D <= "00000000";	-- 0x1983
		when 006532 => D <= "11011101";	-- 0x1984
		when 006533 => D <= "11100001";	-- 0x1985
		when 006534 => D <= "11100101";	-- 0x1986
		when 006535 => D <= "11011101";	-- 0x1987
		when 006536 => D <= "01111110";	-- 0x1988
		when 006537 => D <= "00000000";	-- 0x1989
		when 006538 => D <= "10110111";	-- 0x198A
		when 006539 => D <= "11001010";	-- 0x198B
		when 006540 => D <= "10011010";	-- 0x198C
		when 006541 => D <= "00111001";	-- 0x198D
		when 006542 => D <= "01001111";	-- 0x198E
		when 006543 => D <= "11001101";	-- 0x198F
		when 006544 => D <= "10110111";	-- 0x1990
		when 006545 => D <= "00110000";	-- 0x1991
		when 006546 => D <= "11011101";	-- 0x1992
		when 006547 => D <= "00100011";	-- 0x1993
		when 006548 => D <= "11011101";	-- 0x1994
		when 006549 => D <= "01111110";	-- 0x1995
		when 006550 => D <= "00000000";	-- 0x1996
		when 006551 => D <= "11000011";	-- 0x1997
		when 006552 => D <= "10001010";	-- 0x1998
		when 006553 => D <= "00111001";	-- 0x1999
		when 006554 => D <= "11011101";	-- 0x199A
		when 006555 => D <= "00100011";	-- 0x199B
		when 006556 => D <= "11001101";	-- 0x199C
		when 006557 => D <= "11101111";	-- 0x199D
		when 006558 => D <= "00110000";	-- 0x199E
		when 006559 => D <= "11100001";	-- 0x199F
		when 006560 => D <= "01111101";	-- 0x19A0
		when 006561 => D <= "11111110";	-- 0x19A1
		when 006562 => D <= "10001010";	-- 0x19A2
		when 006563 => D <= "11000010";	-- 0x19A3
		when 006564 => D <= "01110011";	-- 0x19A4
		when 006565 => D <= "00111001";	-- 0x19A5
		when 006566 => D <= "11011101";	-- 0x19A6
		when 006567 => D <= "11100001";	-- 0x19A7
		when 006568 => D <= "11000011";	-- 0x19A8
		when 006569 => D <= "11101100";	-- 0x19A9
		when 006570 => D <= "00111001";	-- 0x19AA
		when 006571 => D <= "00100001";	-- 0x19AB
		when 006572 => D <= "01001111";	-- 0x19AC
		when 006573 => D <= "10000011";	-- 0x19AD
		when 006574 => D <= "11100101";	-- 0x19AE
		when 006575 => D <= "00100001";	-- 0x19AF
		when 006576 => D <= "11101100";	-- 0x19B0
		when 006577 => D <= "00111001";	-- 0x19B1
		when 006578 => D <= "11100011";	-- 0x19B2
		when 006579 => D <= "01111110";	-- 0x19B3
		when 006580 => D <= "10110111";	-- 0x19B4
		when 006581 => D <= "11001000";	-- 0x19B5
		when 006582 => D <= "11001011";	-- 0x19B6
		when 006583 => D <= "01111111";	-- 0x19B7
		when 006584 => D <= "11001010";	-- 0x19B8
		when 006585 => D <= "11100100";	-- 0x19B9
		when 006586 => D <= "00111001";	-- 0x19BA
		when 006587 => D <= "11001011";	-- 0x19BB
		when 006588 => D <= "10111111";	-- 0x19BC
		when 006589 => D <= "01001111";	-- 0x19BD
		when 006590 => D <= "11001101";	-- 0x19BE
		when 006591 => D <= "10110111";	-- 0x19BF
		when 006592 => D <= "00110000";	-- 0x19C0
		when 006593 => D <= "00100011";	-- 0x19C1
		when 006594 => D <= "00100011";	-- 0x19C2
		when 006595 => D <= "00100011";	-- 0x19C3
		when 006596 => D <= "01111110";	-- 0x19C4
		when 006597 => D <= "11111110";	-- 0x19C5
		when 006598 => D <= "00000001";	-- 0x19C6
		when 006599 => D <= "11000010";	-- 0x19C7
		when 006600 => D <= "11010101";	-- 0x19C8
		when 006601 => D <= "00111001";	-- 0x19C9
		when 006602 => D <= "11100101";	-- 0x19CA
		when 006603 => D <= "00100001";	-- 0x19CB
		when 006604 => D <= "11101101";	-- 0x19CC
		when 006605 => D <= "00111001";	-- 0x19CD
		when 006606 => D <= "11001101";	-- 0x19CE
		when 006607 => D <= "10110010";	-- 0x19CF
		when 006608 => D <= "00111110";	-- 0x19D0
		when 006609 => D <= "11100001";	-- 0x19D1
		when 006610 => D <= "11000011";	-- 0x19D2
		when 006611 => D <= "11011101";	-- 0x19D3
		when 006612 => D <= "00111001";	-- 0x19D4
		when 006613 => D <= "11100101";	-- 0x19D5
		when 006614 => D <= "00100001";	-- 0x19D6
		when 006615 => D <= "11111011";	-- 0x19D7
		when 006616 => D <= "00111001";	-- 0x19D8
		when 006617 => D <= "11001101";	-- 0x19D9
		when 006618 => D <= "10110010";	-- 0x19DA
		when 006619 => D <= "00111110";	-- 0x19DB
		when 006620 => D <= "11100001";	-- 0x19DC
		when 006621 => D <= "00100011";	-- 0x19DD
		when 006622 => D <= "11001101";	-- 0x19DE
		when 006623 => D <= "11101111";	-- 0x19DF
		when 006624 => D <= "00110000";	-- 0x19E0
		when 006625 => D <= "11000011";	-- 0x19E1
		when 006626 => D <= "11101001";	-- 0x19E2
		when 006627 => D <= "00111001";	-- 0x19E3
		when 006628 => D <= "01001111";	-- 0x19E4
		when 006629 => D <= "11001101";	-- 0x19E5
		when 006630 => D <= "10110111";	-- 0x19E6
		when 006631 => D <= "00110000";	-- 0x19E7
		when 006632 => D <= "00100011";	-- 0x19E8
		when 006633 => D <= "11000011";	-- 0x19E9
		when 006634 => D <= "10110011";	-- 0x19EA
		when 006635 => D <= "00111001";	-- 0x19EB
		when 006636 => D <= "11001001";	-- 0x19EC
		when 006637 => D <= "00100000";	-- 0x19ED
		when 006638 => D <= "01101001";	-- 0x19EE
		when 006639 => D <= "01110011";	-- 0x19EF
		when 006640 => D <= "01110100";	-- 0x19F0
		when 006641 => D <= "00100000";	-- 0x19F1
		when 006642 => D <= "01010110";	-- 0x19F2
		when 006643 => D <= "01100001";	-- 0x19F3
		when 006644 => D <= "01110010";	-- 0x19F4
		when 006645 => D <= "01101001";	-- 0x19F5
		when 006646 => D <= "01100001";	-- 0x19F6
		when 006647 => D <= "01100010";	-- 0x19F7
		when 006648 => D <= "01101100";	-- 0x19F8
		when 006649 => D <= "01100101";	-- 0x19F9
		when 006650 => D <= "00000000";	-- 0x19FA
		when 006651 => D <= "00100000";	-- 0x19FB
		when 006652 => D <= "01101001";	-- 0x19FC
		when 006653 => D <= "01110011";	-- 0x19FD
		when 006654 => D <= "01110100";	-- 0x19FE
		when 006655 => D <= "00100000";	-- 0x19FF
		when 006656 => D <= "01100111";	-- 0x1A00
		when 006657 => D <= "01100101";	-- 0x1A01
		when 006658 => D <= "01101100";	-- 0x1A02
		when 006659 => D <= "01100101";	-- 0x1A03
		when 006660 => D <= "01110010";	-- 0x1A04
		when 006661 => D <= "01101110";	-- 0x1A05
		when 006662 => D <= "01110100";	-- 0x1A06
		when 006663 => D <= "00000000";	-- 0x1A07
		when 006664 => D <= "00111110";	-- 0x1A08
		when 006665 => D <= "00000001";	-- 0x1A09
		when 006666 => D <= "00011000";	-- 0x1A0A
		when 006667 => D <= "00000001";	-- 0x1A0B
		when 006668 => D <= "10101111";	-- 0x1A0C
		when 006669 => D <= "00110010";	-- 0x1A0D
		when 006670 => D <= "01000000";	-- 0x1A0E
		when 006671 => D <= "10000011";	-- 0x1A0F
		when 006672 => D <= "11001101";	-- 0x1A10
		when 006673 => D <= "11000110";	-- 0x1A11
		when 006674 => D <= "00100000";	-- 0x1A12
		when 006675 => D <= "11111110";	-- 0x1A13
		when 006676 => D <= "11111111";	-- 0x1A14
		when 006677 => D <= "11000010";	-- 0x1A15
		when 006678 => D <= "00010000";	-- 0x1A16
		when 006679 => D <= "00111010";	-- 0x1A17
		when 006680 => D <= "11001101";	-- 0x1A18
		when 006681 => D <= "11000110";	-- 0x1A19
		when 006682 => D <= "00100000";	-- 0x1A1A
		when 006683 => D <= "10110111";	-- 0x1A1B
		when 006684 => D <= "11000010";	-- 0x1A1C
		when 006685 => D <= "00011000";	-- 0x1A1D
		when 006686 => D <= "00111010";	-- 0x1A1E
		when 006687 => D <= "11001101";	-- 0x1A1F
		when 006688 => D <= "11000110";	-- 0x1A20
		when 006689 => D <= "00100000";	-- 0x1A21
		when 006690 => D <= "11111110";	-- 0x1A22
		when 006691 => D <= "00101111";	-- 0x1A23
		when 006692 => D <= "11000010";	-- 0x1A24
		when 006693 => D <= "00010000";	-- 0x1A25
		when 006694 => D <= "00111010";	-- 0x1A26
		when 006695 => D <= "11001101";	-- 0x1A27
		when 006696 => D <= "11000110";	-- 0x1A28
		when 006697 => D <= "00100000";	-- 0x1A29
		when 006698 => D <= "11111110";	-- 0x1A2A
		when 006699 => D <= "00001101";	-- 0x1A2B
		when 006700 => D <= "11001010";	-- 0x1A2C
		when 006701 => D <= "00111001";	-- 0x1A2D
		when 006702 => D <= "00111010";	-- 0x1A2E
		when 006703 => D <= "01001111";	-- 0x1A2F
		when 006704 => D <= "11001101";	-- 0x1A30
		when 006705 => D <= "10110111";	-- 0x1A31
		when 006706 => D <= "00110000";	-- 0x1A32
		when 006707 => D <= "11001101";	-- 0x1A33
		when 006708 => D <= "11000110";	-- 0x1A34
		when 006709 => D <= "00100000";	-- 0x1A35
		when 006710 => D <= "11000011";	-- 0x1A36
		when 006711 => D <= "00101010";	-- 0x1A37
		when 006712 => D <= "00111010";	-- 0x1A38
		when 006713 => D <= "00001110";	-- 0x1A39
		when 006714 => D <= "00111010";	-- 0x1A3A
		when 006715 => D <= "11001101";	-- 0x1A3B
		when 006716 => D <= "01001010";	-- 0x1A3C
		when 006717 => D <= "00111010";	-- 0x1A3D
		when 006718 => D <= "11011010";	-- 0x1A3E
		when 006719 => D <= "01000110";	-- 0x1A3F
		when 006720 => D <= "00111010";	-- 0x1A40
		when 006721 => D <= "00001110";	-- 0x1A41
		when 006722 => D <= "00100100";	-- 0x1A42
		when 006723 => D <= "11001101";	-- 0x1A43
		when 006724 => D <= "01001010";	-- 0x1A44
		when 006725 => D <= "00111010";	-- 0x1A45
		when 006726 => D <= "11001101";	-- 0x1A46
		when 006727 => D <= "10110010";	-- 0x1A47
		when 006728 => D <= "00111110";	-- 0x1A48
		when 006729 => D <= "11001001";	-- 0x1A49
		when 006730 => D <= "11001101";	-- 0x1A4A
		when 006731 => D <= "11000110";	-- 0x1A4B
		when 006732 => D <= "00100000";	-- 0x1A4C
		when 006733 => D <= "10110111";	-- 0x1A4D
		when 006734 => D <= "11000010";	-- 0x1A4E
		when 006735 => D <= "01001010";	-- 0x1A4F
		when 006736 => D <= "00111010";	-- 0x1A50
		when 006737 => D <= "11001101";	-- 0x1A51
		when 006738 => D <= "11000110";	-- 0x1A52
		when 006739 => D <= "00100000";	-- 0x1A53
		when 006740 => D <= "10111001";	-- 0x1A54
		when 006741 => D <= "11000010";	-- 0x1A55
		when 006742 => D <= "01001010";	-- 0x1A56
		when 006743 => D <= "00111010";	-- 0x1A57
		when 006744 => D <= "00100001";	-- 0x1A58
		when 006745 => D <= "00000000";	-- 0x1A59
		when 006746 => D <= "00000000";	-- 0x1A5A
		when 006747 => D <= "11001101";	-- 0x1A5B
		when 006748 => D <= "11000110";	-- 0x1A5C
		when 006749 => D <= "00100000";	-- 0x1A5D
		when 006750 => D <= "01010111";	-- 0x1A5E
		when 006751 => D <= "11001101";	-- 0x1A5F
		when 006752 => D <= "11000110";	-- 0x1A60
		when 006753 => D <= "00100000";	-- 0x1A61
		when 006754 => D <= "01011111";	-- 0x1A62
		when 006755 => D <= "11101101";	-- 0x1A63
		when 006756 => D <= "01010011";	-- 0x1A64
		when 006757 => D <= "11100010";	-- 0x1A65
		when 006758 => D <= "10000010";	-- 0x1A66
		when 006759 => D <= "00011001";	-- 0x1A67
		when 006760 => D <= "11010101";	-- 0x1A68
		when 006761 => D <= "11001101";	-- 0x1A69
		when 006762 => D <= "11000110";	-- 0x1A6A
		when 006763 => D <= "00100000";	-- 0x1A6B
		when 006764 => D <= "01010111";	-- 0x1A6C
		when 006765 => D <= "11001101";	-- 0x1A6D
		when 006766 => D <= "11000110";	-- 0x1A6E
		when 006767 => D <= "00100000";	-- 0x1A6F
		when 006768 => D <= "01011111";	-- 0x1A70
		when 006769 => D <= "11101101";	-- 0x1A71
		when 006770 => D <= "01010011";	-- 0x1A72
		when 006771 => D <= "11100100";	-- 0x1A73
		when 006772 => D <= "10000010";	-- 0x1A74
		when 006773 => D <= "00011001";	-- 0x1A75
		when 006774 => D <= "11010001";	-- 0x1A76
		when 006775 => D <= "11100101";	-- 0x1A77
		when 006776 => D <= "00100001";	-- 0x1A78
		when 006777 => D <= "10100110";	-- 0x1A79
		when 006778 => D <= "00111010";	-- 0x1A7A
		when 006779 => D <= "11100011";	-- 0x1A7B
		when 006780 => D <= "11001101";	-- 0x1A7C
		when 006781 => D <= "11000110";	-- 0x1A7D
		when 006782 => D <= "00100000";	-- 0x1A7E
		when 006783 => D <= "01001111";	-- 0x1A7F
		when 006784 => D <= "00000110";	-- 0x1A80
		when 006785 => D <= "00000000";	-- 0x1A81
		when 006786 => D <= "00001001";	-- 0x1A82
		when 006787 => D <= "00111010";	-- 0x1A83
		when 006788 => D <= "01000000";	-- 0x1A84
		when 006789 => D <= "10000011";	-- 0x1A85
		when 006790 => D <= "10110111";	-- 0x1A86
		when 006791 => D <= "11000010";	-- 0x1A87
		when 006792 => D <= "10001100";	-- 0x1A88
		when 006793 => D <= "00111010";	-- 0x1A89
		when 006794 => D <= "01111001";	-- 0x1A8A
		when 006795 => D <= "00010010";	-- 0x1A8B
		when 006796 => D <= "00011010";	-- 0x1A8C
		when 006797 => D <= "10111001";	-- 0x1A8D
		when 006798 => D <= "11001010";	-- 0x1A8E
		when 006799 => D <= "10010011";	-- 0x1A8F
		when 006800 => D <= "00111010";	-- 0x1A90
		when 006801 => D <= "00110111";	-- 0x1A91
		when 006802 => D <= "11001001";	-- 0x1A92
		when 006803 => D <= "11100101";	-- 0x1A93
		when 006804 => D <= "00101010";	-- 0x1A94
		when 006805 => D <= "11100100";	-- 0x1A95
		when 006806 => D <= "10000010";	-- 0x1A96
		when 006807 => D <= "10101111";	-- 0x1A97
		when 006808 => D <= "11101101";	-- 0x1A98
		when 006809 => D <= "01010010";	-- 0x1A99
		when 006810 => D <= "01111100";	-- 0x1A9A
		when 006811 => D <= "10110101";	-- 0x1A9B
		when 006812 => D <= "11100001";	-- 0x1A9C
		when 006813 => D <= "11000010";	-- 0x1A9D
		when 006814 => D <= "10100010";	-- 0x1A9E
		when 006815 => D <= "00111010";	-- 0x1A9F
		when 006816 => D <= "10101111";	-- 0x1AA0
		when 006817 => D <= "11001001";	-- 0x1AA1
		when 006818 => D <= "00010011";	-- 0x1AA2
		when 006819 => D <= "11000011";	-- 0x1AA3
		when 006820 => D <= "01111100";	-- 0x1AA4
		when 006821 => D <= "00111010";	-- 0x1AA5
		when 006822 => D <= "11101011";	-- 0x1AA6
		when 006823 => D <= "00100001";	-- 0x1AA7
		when 006824 => D <= "11000100";	-- 0x1AA8
		when 006825 => D <= "00111010";	-- 0x1AA9
		when 006826 => D <= "00110000";	-- 0x1AAA
		when 006827 => D <= "00000101";	-- 0x1AAB
		when 006828 => D <= "00100001";	-- 0x1AAC
		when 006829 => D <= "11011000";	-- 0x1AAD
		when 006830 => D <= "00111010";	-- 0x1AAE
		when 006831 => D <= "00110111";	-- 0x1AAF
		when 006832 => D <= "11001001";	-- 0x1AB0
		when 006833 => D <= "11001101";	-- 0x1AB1
		when 006834 => D <= "11000110";	-- 0x1AB2
		when 006835 => D <= "00100000";	-- 0x1AB3
		when 006836 => D <= "10111010";	-- 0x1AB4
		when 006837 => D <= "00101000";	-- 0x1AB5
		when 006838 => D <= "00000101";	-- 0x1AB6
		when 006839 => D <= "00100001";	-- 0x1AB7
		when 006840 => D <= "11001010";	-- 0x1AB8
		when 006841 => D <= "00111010";	-- 0x1AB9
		when 006842 => D <= "00110111";	-- 0x1ABA
		when 006843 => D <= "11001001";	-- 0x1ABB
		when 006844 => D <= "11001101";	-- 0x1ABC
		when 006845 => D <= "11000110";	-- 0x1ABD
		when 006846 => D <= "00100000";	-- 0x1ABE
		when 006847 => D <= "10111011";	-- 0x1ABF
		when 006848 => D <= "00100000";	-- 0x1AC0
		when 006849 => D <= "11110101";	-- 0x1AC1
		when 006850 => D <= "10101111";	-- 0x1AC2
		when 006851 => D <= "11001001";	-- 0x1AC3
		when 006852 => D <= "00100000";	-- 0x1AC4
		when 006853 => D <= "01001111";	-- 0x1AC5
		when 006854 => D <= "01101011";	-- 0x1AC6
		when 006855 => D <= "00001101";	-- 0x1AC7
		when 006856 => D <= "00001010";	-- 0x1AC8
		when 006857 => D <= "00000000";	-- 0x1AC9
		when 006858 => D <= "00100000";	-- 0x1ACA
		when 006859 => D <= "01000110";	-- 0x1ACB
		when 006860 => D <= "01100101";	-- 0x1ACC
		when 006861 => D <= "01101000";	-- 0x1ACD
		when 006862 => D <= "01101100";	-- 0x1ACE
		when 006863 => D <= "01100101";	-- 0x1ACF
		when 006864 => D <= "01110010";	-- 0x1AD0
		when 006865 => D <= "00100000";	-- 0x1AD1
		when 006866 => D <= "01000011";	-- 0x1AD2
		when 006867 => D <= "01000001";	-- 0x1AD3
		when 006868 => D <= "01010011";	-- 0x1AD4
		when 006869 => D <= "00001101";	-- 0x1AD5
		when 006870 => D <= "00001010";	-- 0x1AD6
		when 006871 => D <= "00000000";	-- 0x1AD7
		when 006872 => D <= "00100000";	-- 0x1AD8
		when 006873 => D <= "01000110";	-- 0x1AD9
		when 006874 => D <= "01100101";	-- 0x1ADA
		when 006875 => D <= "01101000";	-- 0x1ADB
		when 006876 => D <= "01101100";	-- 0x1ADC
		when 006877 => D <= "01100101";	-- 0x1ADD
		when 006878 => D <= "01110010";	-- 0x1ADE
		when 006879 => D <= "00100000";	-- 0x1ADF
		when 006880 => D <= "01010110";	-- 0x1AE0
		when 006881 => D <= "01100111";	-- 0x1AE1
		when 006882 => D <= "01101100";	-- 0x1AE2
		when 006883 => D <= "00001101";	-- 0x1AE3
		when 006884 => D <= "00001010";	-- 0x1AE4
		when 006885 => D <= "00000000";	-- 0x1AE5
		when 006886 => D <= "00000110";	-- 0x1AE6
		when 006887 => D <= "00101000";	-- 0x1AE7
		when 006888 => D <= "00001110";	-- 0x1AE8
		when 006889 => D <= "11111111";	-- 0x1AE9
		when 006890 => D <= "11001101";	-- 0x1AEA
		when 006891 => D <= "11001111";	-- 0x1AEB
		when 006892 => D <= "00100000";	-- 0x1AEC
		when 006893 => D <= "00000101";	-- 0x1AED
		when 006894 => D <= "11000010";	-- 0x1AEE
		when 006895 => D <= "11101000";	-- 0x1AEF
		when 006896 => D <= "00111010";	-- 0x1AF0
		when 006897 => D <= "00001110";	-- 0x1AF1
		when 006898 => D <= "00000000";	-- 0x1AF2
		when 006899 => D <= "11001101";	-- 0x1AF3
		when 006900 => D <= "11001111";	-- 0x1AF4
		when 006901 => D <= "00100000";	-- 0x1AF5
		when 006902 => D <= "00001110";	-- 0x1AF6
		when 006903 => D <= "00101111";	-- 0x1AF7
		when 006904 => D <= "11001101";	-- 0x1AF8
		when 006905 => D <= "11001111";	-- 0x1AF9
		when 006906 => D <= "00100000";	-- 0x1AFA
		when 006907 => D <= "11011101";	-- 0x1AFB
		when 006908 => D <= "01111110";	-- 0x1AFC
		when 006909 => D <= "00000000";	-- 0x1AFD
		when 006910 => D <= "10110111";	-- 0x1AFE
		when 006911 => D <= "11001010";	-- 0x1AFF
		when 006912 => D <= "00001101";	-- 0x1B00
		when 006913 => D <= "00111011";	-- 0x1B01
		when 006914 => D <= "11011101";	-- 0x1B02
		when 006915 => D <= "01001110";	-- 0x1B03
		when 006916 => D <= "00000000";	-- 0x1B04
		when 006917 => D <= "11001101";	-- 0x1B05
		when 006918 => D <= "11001111";	-- 0x1B06
		when 006919 => D <= "00100000";	-- 0x1B07
		when 006920 => D <= "11011101";	-- 0x1B08
		when 006921 => D <= "00100011";	-- 0x1B09
		when 006922 => D <= "11000011";	-- 0x1B0A
		when 006923 => D <= "11111011";	-- 0x1B0B
		when 006924 => D <= "00111010";	-- 0x1B0C
		when 006925 => D <= "00001110";	-- 0x1B0D
		when 006926 => D <= "00001101";	-- 0x1B0E
		when 006927 => D <= "11001101";	-- 0x1B0F
		when 006928 => D <= "11001111";	-- 0x1B10
		when 006929 => D <= "00100000";	-- 0x1B11
		when 006930 => D <= "00001110";	-- 0x1B12
		when 006931 => D <= "00111010";	-- 0x1B13
		when 006932 => D <= "00101010";	-- 0x1B14
		when 006933 => D <= "01000001";	-- 0x1B15
		when 006934 => D <= "10000011";	-- 0x1B16
		when 006935 => D <= "00100010";	-- 0x1B17
		when 006936 => D <= "11100010";	-- 0x1B18
		when 006937 => D <= "10000010";	-- 0x1B19
		when 006938 => D <= "00101010";	-- 0x1B1A
		when 006939 => D <= "01000011";	-- 0x1B1B
		when 006940 => D <= "10000011";	-- 0x1B1C
		when 006941 => D <= "00100010";	-- 0x1B1D
		when 006942 => D <= "11100100";	-- 0x1B1E
		when 006943 => D <= "10000010";	-- 0x1B1F
		when 006944 => D <= "11001101";	-- 0x1B20
		when 006945 => D <= "01000000";	-- 0x1B21
		when 006946 => D <= "00111011";	-- 0x1B22
		when 006947 => D <= "00001110";	-- 0x1B23
		when 006948 => D <= "00100100";	-- 0x1B24
		when 006949 => D <= "00100001";	-- 0x1B25
		when 006950 => D <= "01000001";	-- 0x1B26
		when 006951 => D <= "10000011";	-- 0x1B27
		when 006952 => D <= "00100010";	-- 0x1B28
		when 006953 => D <= "11100010";	-- 0x1B29
		when 006954 => D <= "10000010";	-- 0x1B2A
		when 006955 => D <= "00101010";	-- 0x1B2B
		when 006956 => D <= "01001001";	-- 0x1B2C
		when 006957 => D <= "10000011";	-- 0x1B2D
		when 006958 => D <= "00100010";	-- 0x1B2E
		when 006959 => D <= "11100100";	-- 0x1B2F
		when 006960 => D <= "10000010";	-- 0x1B30
		when 006961 => D <= "11001101";	-- 0x1B31
		when 006962 => D <= "01000000";	-- 0x1B32
		when 006963 => D <= "00111011";	-- 0x1B33
		when 006964 => D <= "00000110";	-- 0x1B34
		when 006965 => D <= "00010100";	-- 0x1B35
		when 006966 => D <= "00001110";	-- 0x1B36
		when 006967 => D <= "11111111";	-- 0x1B37
		when 006968 => D <= "11001101";	-- 0x1B38
		when 006969 => D <= "11001111";	-- 0x1B39
		when 006970 => D <= "00100000";	-- 0x1B3A
		when 006971 => D <= "00000101";	-- 0x1B3B
		when 006972 => D <= "11000010";	-- 0x1B3C
		when 006973 => D <= "00110110";	-- 0x1B3D
		when 006974 => D <= "00111011";	-- 0x1B3E
		when 006975 => D <= "11001001";	-- 0x1B3F
		when 006976 => D <= "11000101";	-- 0x1B40
		when 006977 => D <= "00000110";	-- 0x1B41
		when 006978 => D <= "00010100";	-- 0x1B42
		when 006979 => D <= "00001110";	-- 0x1B43
		when 006980 => D <= "11111111";	-- 0x1B44
		when 006981 => D <= "11001101";	-- 0x1B45
		when 006982 => D <= "11001111";	-- 0x1B46
		when 006983 => D <= "00100000";	-- 0x1B47
		when 006984 => D <= "00000101";	-- 0x1B48
		when 006985 => D <= "11000010";	-- 0x1B49
		when 006986 => D <= "01000011";	-- 0x1B4A
		when 006987 => D <= "00111011";	-- 0x1B4B
		when 006988 => D <= "00001110";	-- 0x1B4C
		when 006989 => D <= "00000000";	-- 0x1B4D
		when 006990 => D <= "11001101";	-- 0x1B4E
		when 006991 => D <= "11001111";	-- 0x1B4F
		when 006992 => D <= "00100000";	-- 0x1B50
		when 006993 => D <= "11000001";	-- 0x1B51
		when 006994 => D <= "11001101";	-- 0x1B52
		when 006995 => D <= "11001111";	-- 0x1B53
		when 006996 => D <= "00100000";	-- 0x1B54
		when 006997 => D <= "00100001";	-- 0x1B55
		when 006998 => D <= "00000000";	-- 0x1B56
		when 006999 => D <= "00000000";	-- 0x1B57
		when 007000 => D <= "11101101";	-- 0x1B58
		when 007001 => D <= "01011011";	-- 0x1B59
		when 007002 => D <= "11100010";	-- 0x1B5A
		when 007003 => D <= "10000010";	-- 0x1B5B
		when 007004 => D <= "00011001";	-- 0x1B5C
		when 007005 => D <= "11010101";	-- 0x1B5D
		when 007006 => D <= "01001010";	-- 0x1B5E
		when 007007 => D <= "11001101";	-- 0x1B5F
		when 007008 => D <= "11001111";	-- 0x1B60
		when 007009 => D <= "00100000";	-- 0x1B61
		when 007010 => D <= "01001011";	-- 0x1B62
		when 007011 => D <= "11001101";	-- 0x1B63
		when 007012 => D <= "11001111";	-- 0x1B64
		when 007013 => D <= "00100000";	-- 0x1B65
		when 007014 => D <= "11101101";	-- 0x1B66
		when 007015 => D <= "01011011";	-- 0x1B67
		when 007016 => D <= "11100100";	-- 0x1B68
		when 007017 => D <= "10000010";	-- 0x1B69
		when 007018 => D <= "00011001";	-- 0x1B6A
		when 007019 => D <= "01001010";	-- 0x1B6B
		when 007020 => D <= "11001101";	-- 0x1B6C
		when 007021 => D <= "11001111";	-- 0x1B6D
		when 007022 => D <= "00100000";	-- 0x1B6E
		when 007023 => D <= "01001011";	-- 0x1B6F
		when 007024 => D <= "11001101";	-- 0x1B70
		when 007025 => D <= "11001111";	-- 0x1B71
		when 007026 => D <= "00100000";	-- 0x1B72
		when 007027 => D <= "11010001";	-- 0x1B73
		when 007028 => D <= "11100101";	-- 0x1B74
		when 007029 => D <= "00100001";	-- 0x1B75
		when 007030 => D <= "10010000";	-- 0x1B76
		when 007031 => D <= "00111011";	-- 0x1B77
		when 007032 => D <= "11100011";	-- 0x1B78
		when 007033 => D <= "00011010";	-- 0x1B79
		when 007034 => D <= "01001111";	-- 0x1B7A
		when 007035 => D <= "00000110";	-- 0x1B7B
		when 007036 => D <= "00000000";	-- 0x1B7C
		when 007037 => D <= "00001001";	-- 0x1B7D
		when 007038 => D <= "11001101";	-- 0x1B7E
		when 007039 => D <= "11001111";	-- 0x1B7F
		when 007040 => D <= "00100000";	-- 0x1B80
		when 007041 => D <= "11100101";	-- 0x1B81
		when 007042 => D <= "00101010";	-- 0x1B82
		when 007043 => D <= "11100100";	-- 0x1B83
		when 007044 => D <= "10000010";	-- 0x1B84
		when 007045 => D <= "10101111";	-- 0x1B85
		when 007046 => D <= "11101101";	-- 0x1B86
		when 007047 => D <= "01010010";	-- 0x1B87
		when 007048 => D <= "01111100";	-- 0x1B88
		when 007049 => D <= "10110101";	-- 0x1B89
		when 007050 => D <= "11100001";	-- 0x1B8A
		when 007051 => D <= "11001000";	-- 0x1B8B
		when 007052 => D <= "00010011";	-- 0x1B8C
		when 007053 => D <= "11000011";	-- 0x1B8D
		when 007054 => D <= "01111001";	-- 0x1B8E
		when 007055 => D <= "00111011";	-- 0x1B8F
		when 007056 => D <= "01001100";	-- 0x1B90
		when 007057 => D <= "11001101";	-- 0x1B91
		when 007058 => D <= "11001111";	-- 0x1B92
		when 007059 => D <= "00100000";	-- 0x1B93
		when 007060 => D <= "01001101";	-- 0x1B94
		when 007061 => D <= "11001101";	-- 0x1B95
		when 007062 => D <= "11001111";	-- 0x1B96
		when 007063 => D <= "00100000";	-- 0x1B97
		when 007064 => D <= "11001001";	-- 0x1B98
		when 007065 => D <= "11001101";	-- 0x1B99
		when 007066 => D <= "11001100";	-- 0x1B9A
		when 007067 => D <= "00100111";	-- 0x1B9B
		when 007068 => D <= "11011101";	-- 0x1B9C
		when 007069 => D <= "01111110";	-- 0x1B9D
		when 007070 => D <= "00000000";	-- 0x1B9E
		when 007071 => D <= "11111110";	-- 0x1B9F
		when 007072 => D <= "00100010";	-- 0x1BA0
		when 007073 => D <= "11001010";	-- 0x1BA1
		when 007074 => D <= "10100110";	-- 0x1BA2
		when 007075 => D <= "00111011";	-- 0x1BA3
		when 007076 => D <= "00110111";	-- 0x1BA4
		when 007077 => D <= "11001001";	-- 0x1BA5
		when 007078 => D <= "11011101";	-- 0x1BA6
		when 007079 => D <= "00100011";	-- 0x1BA7
		when 007080 => D <= "11011101";	-- 0x1BA8
		when 007081 => D <= "11100101";	-- 0x1BA9
		when 007082 => D <= "11011101";	-- 0x1BAA
		when 007083 => D <= "01111110";	-- 0x1BAB
		when 007084 => D <= "00000000";	-- 0x1BAC
		when 007085 => D <= "11111110";	-- 0x1BAD
		when 007086 => D <= "01111011";	-- 0x1BAE
		when 007087 => D <= "00110000";	-- 0x1BAF
		when 007088 => D <= "00000101";	-- 0x1BB0
		when 007089 => D <= "11111110";	-- 0x1BB1
		when 007090 => D <= "01100001";	-- 0x1BB2
		when 007091 => D <= "11010010";	-- 0x1BB3
		when 007092 => D <= "11000000";	-- 0x1BB4
		when 007093 => D <= "00111011";	-- 0x1BB5
		when 007094 => D <= "11111110";	-- 0x1BB6
		when 007095 => D <= "01011011";	-- 0x1BB7
		when 007096 => D <= "11010010";	-- 0x1BB8
		when 007097 => D <= "11111000";	-- 0x1BB9
		when 007098 => D <= "00111011";	-- 0x1BBA
		when 007099 => D <= "11111110";	-- 0x1BBB
		when 007100 => D <= "01000001";	-- 0x1BBC
		when 007101 => D <= "11011010";	-- 0x1BBD
		when 007102 => D <= "11111000";	-- 0x1BBE
		when 007103 => D <= "00111011";	-- 0x1BBF
		when 007104 => D <= "10101111";	-- 0x1BC0
		when 007105 => D <= "11011010";	-- 0x1BC1
		when 007106 => D <= "11001111";	-- 0x1BC2
		when 007107 => D <= "00111011";	-- 0x1BC3
		when 007108 => D <= "11011101";	-- 0x1BC4
		when 007109 => D <= "00100011";	-- 0x1BC5
		when 007110 => D <= "11011101";	-- 0x1BC6
		when 007111 => D <= "01111110";	-- 0x1BC7
		when 007112 => D <= "00000000";	-- 0x1BC8
		when 007113 => D <= "11001101";	-- 0x1BC9
		when 007114 => D <= "10111100";	-- 0x1BCA
		when 007115 => D <= "00101010";	-- 0x1BCB
		when 007116 => D <= "11000011";	-- 0x1BCC
		when 007117 => D <= "11000001";	-- 0x1BCD
		when 007118 => D <= "00111011";	-- 0x1BCE
		when 007119 => D <= "11001101";	-- 0x1BCF
		when 007120 => D <= "00100010";	-- 0x1BD0
		when 007121 => D <= "00111100";	-- 0x1BD1
		when 007122 => D <= "11011010";	-- 0x1BD2
		when 007123 => D <= "11110010";	-- 0x1BD3
		when 007124 => D <= "00111011";	-- 0x1BD4
		when 007125 => D <= "11011101";	-- 0x1BD5
		when 007126 => D <= "11100011";	-- 0x1BD6
		when 007127 => D <= "00111110";	-- 0x1BD7
		when 007128 => D <= "00000001";	-- 0x1BD8
		when 007129 => D <= "11100101";	-- 0x1BD9
		when 007130 => D <= "11001101";	-- 0x1BDA
		when 007131 => D <= "01110010";	-- 0x1BDB
		when 007132 => D <= "00101011";	-- 0x1BDC
		when 007133 => D <= "11100001";	-- 0x1BDD
		when 007134 => D <= "11010010";	-- 0x1BDE
		when 007135 => D <= "11101011";	-- 0x1BDF
		when 007136 => D <= "00111011";	-- 0x1BE0
		when 007137 => D <= "11111101";	-- 0x1BE1
		when 007138 => D <= "01110101";	-- 0x1BE2
		when 007139 => D <= "00000000";	-- 0x1BE3
		when 007140 => D <= "11111101";	-- 0x1BE4
		when 007141 => D <= "01110100";	-- 0x1BE5
		when 007142 => D <= "00000001";	-- 0x1BE6
		when 007143 => D <= "11111101";	-- 0x1BE7
		when 007144 => D <= "00110110";	-- 0x1BE8
		when 007145 => D <= "00000010";	-- 0x1BE9
		when 007146 => D <= "00000001";	-- 0x1BEA
		when 007147 => D <= "11011101";	-- 0x1BEB
		when 007148 => D <= "11100001";	-- 0x1BEC
		when 007149 => D <= "10101111";	-- 0x1BED
		when 007150 => D <= "11001001";	-- 0x1BEE
		when 007151 => D <= "11000011";	-- 0x1BEF
		when 007152 => D <= "11110101";	-- 0x1BF0
		when 007153 => D <= "00111011";	-- 0x1BF1
		when 007154 => D <= "11000011";	-- 0x1BF2
		when 007155 => D <= "01101110";	-- 0x1BF3
		when 007156 => D <= "00111111";	-- 0x1BF4
		when 007157 => D <= "11000011";	-- 0x1BF5
		when 007158 => D <= "11111000";	-- 0x1BF6
		when 007159 => D <= "00111011";	-- 0x1BF7
		when 007160 => D <= "11011101";	-- 0x1BF8
		when 007161 => D <= "11100001";	-- 0x1BF9
		when 007162 => D <= "00110111";	-- 0x1BFA
		when 007163 => D <= "11001001";	-- 0x1BFB
		when 007164 => D <= "11001101";	-- 0x1BFC
		when 007165 => D <= "00100010";	-- 0x1BFD
		when 007166 => D <= "00111100";	-- 0x1BFE
		when 007167 => D <= "11011010";	-- 0x1BFF
		when 007168 => D <= "01101110";	-- 0x1C00
		when 007169 => D <= "00111111";	-- 0x1C01
		when 007170 => D <= "00010001";	-- 0x1C02
		when 007171 => D <= "00000111";	-- 0x1C03
		when 007172 => D <= "00111100";	-- 0x1C04
		when 007173 => D <= "11010101";	-- 0x1C05
		when 007174 => D <= "11101001";	-- 0x1C06
		when 007175 => D <= "11001001";	-- 0x1C07
		when 007176 => D <= "11000011";	-- 0x1C08
		when 007177 => D <= "01110100";	-- 0x1C09
		when 007178 => D <= "00100010";	-- 0x1C0A
		when 007179 => D <= "11001101";	-- 0x1C0B
		when 007180 => D <= "00100010";	-- 0x1C0C
		when 007181 => D <= "00111100";	-- 0x1C0D
		when 007182 => D <= "11011010";	-- 0x1C0E
		when 007183 => D <= "01101110";	-- 0x1C0F
		when 007184 => D <= "00111111";	-- 0x1C10
		when 007185 => D <= "11100101";	-- 0x1C11
		when 007186 => D <= "11001101";	-- 0x1C12
		when 007187 => D <= "00100010";	-- 0x1C13
		when 007188 => D <= "00111100";	-- 0x1C14
		when 007189 => D <= "11011010";	-- 0x1C15
		when 007190 => D <= "01101110";	-- 0x1C16
		when 007191 => D <= "00111111";	-- 0x1C17
		when 007192 => D <= "11010001";	-- 0x1C18
		when 007193 => D <= "01111101";	-- 0x1C19
		when 007194 => D <= "00110010";	-- 0x1C1A
		when 007195 => D <= "01001001";	-- 0x1C1B
		when 007196 => D <= "10000000";	-- 0x1C1C
		when 007197 => D <= "01111011";	-- 0x1C1D
		when 007198 => D <= "00110010";	-- 0x1C1E
		when 007199 => D <= "01001000";	-- 0x1C1F
		when 007200 => D <= "10000000";	-- 0x1C20
		when 007201 => D <= "11001001";	-- 0x1C21
		when 007202 => D <= "11001101";	-- 0x1C22
		when 007203 => D <= "11001100";	-- 0x1C23
		when 007204 => D <= "00100111";	-- 0x1C24
		when 007205 => D <= "11000011";	-- 0x1C25
		when 007206 => D <= "11111110";	-- 0x1C26
		when 007207 => D <= "00100101";	-- 0x1C27
		when 007208 => D <= "00101010";	-- 0x1C28
		when 007209 => D <= "01000011";	-- 0x1C29
		when 007210 => D <= "10000011";	-- 0x1C2A
		when 007211 => D <= "00010001";	-- 0x1C2B
		when 007212 => D <= "00101000";	-- 0x1C2C
		when 007213 => D <= "00000000";	-- 0x1C2D
		when 007214 => D <= "00011001";	-- 0x1C2E
		when 007215 => D <= "11101011";	-- 0x1C2F
		when 007216 => D <= "00100001";	-- 0x1C30
		when 007217 => D <= "00000000";	-- 0x1C31
		when 007218 => D <= "00000000";	-- 0x1C32
		when 007219 => D <= "00111001";	-- 0x1C33
		when 007220 => D <= "10101111";	-- 0x1C34
		when 007221 => D <= "11101101";	-- 0x1C35
		when 007222 => D <= "01010010";	-- 0x1C36
		when 007223 => D <= "11011010";	-- 0x1C37
		when 007224 => D <= "10000101";	-- 0x1C38
		when 007225 => D <= "00111111";	-- 0x1C39
		when 007226 => D <= "11001001";	-- 0x1C3A
		when 007227 => D <= "11001101";	-- 0x1C3B
		when 007228 => D <= "00101000";	-- 0x1C3C
		when 007229 => D <= "00111100";	-- 0x1C3D
		when 007230 => D <= "11001101";	-- 0x1C3E
		when 007231 => D <= "10001001";	-- 0x1C3F
		when 007232 => D <= "00110000";	-- 0x1C40
		when 007233 => D <= "11001101";	-- 0x1C41
		when 007234 => D <= "11001100";	-- 0x1C42
		when 007235 => D <= "00100111";	-- 0x1C43
		when 007236 => D <= "11111101";	-- 0x1C44
		when 007237 => D <= "00100001";	-- 0x1C45
		when 007238 => D <= "01001111";	-- 0x1C46
		when 007239 => D <= "10000011";	-- 0x1C47
		when 007240 => D <= "11001101";	-- 0x1C48
		when 007241 => D <= "00110101";	-- 0x1C49
		when 007242 => D <= "00101010";	-- 0x1C4A
		when 007243 => D <= "11011010";	-- 0x1C4B
		when 007244 => D <= "11100010";	-- 0x1C4C
		when 007245 => D <= "00111101";	-- 0x1C4D
		when 007246 => D <= "11111110";	-- 0x1C4E
		when 007247 => D <= "00000010";	-- 0x1C4F
		when 007248 => D <= "11000010";	-- 0x1C50
		when 007249 => D <= "11011100";	-- 0x1C51
		when 007250 => D <= "00111101";	-- 0x1C52
		when 007251 => D <= "00111010";	-- 0x1C53
		when 007252 => D <= "00000010";	-- 0x1C54
		when 007253 => D <= "10000000";	-- 0x1C55
		when 007254 => D <= "01000111";	-- 0x1C56
		when 007255 => D <= "00111010";	-- 0x1C57
		when 007256 => D <= "00000011";	-- 0x1C58
		when 007257 => D <= "10000000";	-- 0x1C59
		when 007258 => D <= "01001111";	-- 0x1C5A
		when 007259 => D <= "11000101";	-- 0x1C5B
		when 007260 => D <= "11011101";	-- 0x1C5C
		when 007261 => D <= "00100010";	-- 0x1C5D
		when 007262 => D <= "00001101";	-- 0x1C5E
		when 007263 => D <= "10000000";	-- 0x1C5F
		when 007264 => D <= "00100010";	-- 0x1C60
		when 007265 => D <= "00001111";	-- 0x1C61
		when 007266 => D <= "10000000";	-- 0x1C62
		when 007267 => D <= "11011101";	-- 0x1C63
		when 007268 => D <= "00101010";	-- 0x1C64
		when 007269 => D <= "00001111";	-- 0x1C65
		when 007270 => D <= "10000000";	-- 0x1C66
		when 007271 => D <= "11011101";	-- 0x1C67
		when 007272 => D <= "01111110";	-- 0x1C68
		when 007273 => D <= "00000000";	-- 0x1C69
		when 007274 => D <= "10110111";	-- 0x1C6A
		when 007275 => D <= "11001010";	-- 0x1C6B
		when 007276 => D <= "01111011";	-- 0x1C6C
		when 007277 => D <= "00111100";	-- 0x1C6D
		when 007278 => D <= "11111110";	-- 0x1C6E
		when 007279 => D <= "00111010";	-- 0x1C6F
		when 007280 => D <= "11001010";	-- 0x1C70
		when 007281 => D <= "01111011";	-- 0x1C71
		when 007282 => D <= "00111100";	-- 0x1C72
		when 007283 => D <= "11011101";	-- 0x1C73
		when 007284 => D <= "00100011";	-- 0x1C74
		when 007285 => D <= "11011101";	-- 0x1C75
		when 007286 => D <= "01111110";	-- 0x1C76
		when 007287 => D <= "00000000";	-- 0x1C77
		when 007288 => D <= "11000011";	-- 0x1C78
		when 007289 => D <= "01101010";	-- 0x1C79
		when 007290 => D <= "00111100";	-- 0x1C7A
		when 007291 => D <= "10101111";	-- 0x1C7B
		when 007292 => D <= "00110010";	-- 0x1C7C
		when 007293 => D <= "00010001";	-- 0x1C7D
		when 007294 => D <= "10000000";	-- 0x1C7E
		when 007295 => D <= "11011101";	-- 0x1C7F
		when 007296 => D <= "01111110";	-- 0x1C80
		when 007297 => D <= "00000000";	-- 0x1C81
		when 007298 => D <= "11111110";	-- 0x1C82
		when 007299 => D <= "00111010";	-- 0x1C83
		when 007300 => D <= "11000010";	-- 0x1C84
		when 007301 => D <= "11100010";	-- 0x1C85
		when 007302 => D <= "00111100";	-- 0x1C86
		when 007303 => D <= "11011101";	-- 0x1C87
		when 007304 => D <= "00100011";	-- 0x1C88
		when 007305 => D <= "11011101";	-- 0x1C89
		when 007306 => D <= "00100010";	-- 0x1C8A
		when 007307 => D <= "00001111";	-- 0x1C8B
		when 007308 => D <= "10000000";	-- 0x1C8C
		when 007309 => D <= "11011101";	-- 0x1C8D
		when 007310 => D <= "00101010";	-- 0x1C8E
		when 007311 => D <= "00001101";	-- 0x1C8F
		when 007312 => D <= "10000000";	-- 0x1C90
		when 007313 => D <= "11001101";	-- 0x1C91
		when 007314 => D <= "00100010";	-- 0x1C92
		when 007315 => D <= "00111100";	-- 0x1C93
		when 007316 => D <= "11011010";	-- 0x1C94
		when 007317 => D <= "01101110";	-- 0x1C95
		when 007318 => D <= "00111111";	-- 0x1C96
		when 007319 => D <= "11011101";	-- 0x1C97
		when 007320 => D <= "00100010";	-- 0x1C98
		when 007321 => D <= "00001101";	-- 0x1C99
		when 007322 => D <= "10000000";	-- 0x1C9A
		when 007323 => D <= "00100010";	-- 0x1C9B
		when 007324 => D <= "00010010";	-- 0x1C9C
		when 007325 => D <= "10000000";	-- 0x1C9D
		when 007326 => D <= "11011101";	-- 0x1C9E
		when 007327 => D <= "00101010";	-- 0x1C9F
		when 007328 => D <= "00001111";	-- 0x1CA0
		when 007329 => D <= "10000000";	-- 0x1CA1
		when 007330 => D <= "11011101";	-- 0x1CA2
		when 007331 => D <= "01111110";	-- 0x1CA3
		when 007332 => D <= "00000000";	-- 0x1CA4
		when 007333 => D <= "11001101";	-- 0x1CA5
		when 007334 => D <= "10111100";	-- 0x1CA6
		when 007335 => D <= "00101010";	-- 0x1CA7
		when 007336 => D <= "11011010";	-- 0x1CA8
		when 007337 => D <= "01101110";	-- 0x1CA9
		when 007338 => D <= "00111111";	-- 0x1CAA
		when 007339 => D <= "00111110";	-- 0x1CAB
		when 007340 => D <= "00000001";	-- 0x1CAC
		when 007341 => D <= "11001101";	-- 0x1CAD
		when 007342 => D <= "01110010";	-- 0x1CAE
		when 007343 => D <= "00101011";	-- 0x1CAF
		when 007344 => D <= "11011101";	-- 0x1CB0
		when 007345 => D <= "00100010";	-- 0x1CB1
		when 007346 => D <= "00001111";	-- 0x1CB2
		when 007347 => D <= "10000000";	-- 0x1CB3
		when 007348 => D <= "11010010";	-- 0x1CB4
		when 007349 => D <= "11010101";	-- 0x1CB5
		when 007350 => D <= "00111100";	-- 0x1CB6
		when 007351 => D <= "11111110";	-- 0x1CB7
		when 007352 => D <= "00000010";	-- 0x1CB8
		when 007353 => D <= "11000010";	-- 0x1CB9
		when 007354 => D <= "10111111";	-- 0x1CBA
		when 007355 => D <= "00111100";	-- 0x1CBB
		when 007356 => D <= "11000011";	-- 0x1CBC
		when 007357 => D <= "01101110";	-- 0x1CBD
		when 007358 => D <= "00111111";	-- 0x1CBE
		when 007359 => D <= "11100101";	-- 0x1CBF
		when 007360 => D <= "11111101";	-- 0x1CC0
		when 007361 => D <= "11100101";	-- 0x1CC1
		when 007362 => D <= "11001101";	-- 0x1CC2
		when 007363 => D <= "00101000";	-- 0x1CC3
		when 007364 => D <= "00111100";	-- 0x1CC4
		when 007365 => D <= "00111010";	-- 0x1CC5
		when 007366 => D <= "00010001";	-- 0x1CC6
		when 007367 => D <= "10000000";	-- 0x1CC7
		when 007368 => D <= "00111100";	-- 0x1CC8
		when 007369 => D <= "00110010";	-- 0x1CC9
		when 007370 => D <= "00010001";	-- 0x1CCA
		when 007371 => D <= "10000000";	-- 0x1CCB
		when 007372 => D <= "00101010";	-- 0x1CCC
		when 007373 => D <= "00010010";	-- 0x1CCD
		when 007374 => D <= "10000000";	-- 0x1CCE
		when 007375 => D <= "11111101";	-- 0x1CCF
		when 007376 => D <= "01110101";	-- 0x1CD0
		when 007377 => D <= "00000000";	-- 0x1CD1
		when 007378 => D <= "11111101";	-- 0x1CD2
		when 007379 => D <= "01110100";	-- 0x1CD3
		when 007380 => D <= "00000001";	-- 0x1CD4
		when 007381 => D <= "11011101";	-- 0x1CD5
		when 007382 => D <= "00101010";	-- 0x1CD6
		when 007383 => D <= "00001111";	-- 0x1CD7
		when 007384 => D <= "10000000";	-- 0x1CD8
		when 007385 => D <= "11001101";	-- 0x1CD9
		when 007386 => D <= "11001100";	-- 0x1CDA
		when 007387 => D <= "00100111";	-- 0x1CDB
		when 007388 => D <= "11011101";	-- 0x1CDC
		when 007389 => D <= "01111110";	-- 0x1CDD
		when 007390 => D <= "00000000";	-- 0x1CDE
		when 007391 => D <= "11000011";	-- 0x1CDF
		when 007392 => D <= "10000010";	-- 0x1CE0
		when 007393 => D <= "00111100";	-- 0x1CE1
		when 007394 => D <= "00111010";	-- 0x1CE2
		when 007395 => D <= "00010001";	-- 0x1CE3
		when 007396 => D <= "10000000";	-- 0x1CE4
		when 007397 => D <= "11110101";	-- 0x1CE5
		when 007398 => D <= "11011101";	-- 0x1CE6
		when 007399 => D <= "00101010";	-- 0x1CE7
		when 007400 => D <= "00001101";	-- 0x1CE8
		when 007401 => D <= "10000000";	-- 0x1CE9
		when 007402 => D <= "11011101";	-- 0x1CEA
		when 007403 => D <= "11100101";	-- 0x1CEB
		when 007404 => D <= "11011101";	-- 0x1CEC
		when 007405 => D <= "00101010";	-- 0x1CED
		when 007406 => D <= "00001111";	-- 0x1CEE
		when 007407 => D <= "10000000";	-- 0x1CEF
		when 007408 => D <= "11011101";	-- 0x1CF0
		when 007409 => D <= "01111110";	-- 0x1CF1
		when 007410 => D <= "00000000";	-- 0x1CF2
		when 007411 => D <= "11011101";	-- 0x1CF3
		when 007412 => D <= "00100011";	-- 0x1CF4
		when 007413 => D <= "10110111";	-- 0x1CF5
		when 007414 => D <= "11000010";	-- 0x1CF6
		when 007415 => D <= "11110000";	-- 0x1CF7
		when 007416 => D <= "00111100";	-- 0x1CF8
		when 007417 => D <= "00111110";	-- 0x1CF9
		when 007418 => D <= "11111111";	-- 0x1CFA
		when 007419 => D <= "00110010";	-- 0x1CFB
		when 007420 => D <= "00000010";	-- 0x1CFC
		when 007421 => D <= "10000000";	-- 0x1CFD
		when 007422 => D <= "11011101";	-- 0x1CFE
		when 007423 => D <= "11001011";	-- 0x1CFF
		when 007424 => D <= "00000000";	-- 0x1D00
		when 007425 => D <= "01111110";	-- 0x1D01
		when 007426 => D <= "11001010";	-- 0x1D02
		when 007427 => D <= "10010110";	-- 0x1D03
		when 007428 => D <= "00111101";	-- 0x1D04
		when 007429 => D <= "11111101";	-- 0x1D05
		when 007430 => D <= "00100001";	-- 0x1D06
		when 007431 => D <= "01001111";	-- 0x1D07
		when 007432 => D <= "10000011";	-- 0x1D08
		when 007433 => D <= "11001101";	-- 0x1D09
		when 007434 => D <= "00110101";	-- 0x1D0A
		when 007435 => D <= "00101010";	-- 0x1D0B
		when 007436 => D <= "11011010";	-- 0x1D0C
		when 007437 => D <= "01101110";	-- 0x1D0D
		when 007438 => D <= "00111111";	-- 0x1D0E
		when 007439 => D <= "11111110";	-- 0x1D0F
		when 007440 => D <= "00000010";	-- 0x1D10
		when 007441 => D <= "11000010";	-- 0x1D11
		when 007442 => D <= "01101110";	-- 0x1D12
		when 007443 => D <= "00111111";	-- 0x1D13
		when 007444 => D <= "11011101";	-- 0x1D14
		when 007445 => D <= "00100010";	-- 0x1D15
		when 007446 => D <= "00001101";	-- 0x1D16
		when 007447 => D <= "10000000";	-- 0x1D17
		when 007448 => D <= "00100010";	-- 0x1D18
		when 007449 => D <= "00001111";	-- 0x1D19
		when 007450 => D <= "10000000";	-- 0x1D1A
		when 007451 => D <= "11011101";	-- 0x1D1B
		when 007452 => D <= "00101010";	-- 0x1D1C
		when 007453 => D <= "00001111";	-- 0x1D1D
		when 007454 => D <= "10000000";	-- 0x1D1E
		when 007455 => D <= "11011101";	-- 0x1D1F
		when 007456 => D <= "01111110";	-- 0x1D20
		when 007457 => D <= "00000000";	-- 0x1D21
		when 007458 => D <= "10110111";	-- 0x1D22
		when 007459 => D <= "11001010";	-- 0x1D23
		when 007460 => D <= "00110011";	-- 0x1D24
		when 007461 => D <= "00111101";	-- 0x1D25
		when 007462 => D <= "11111110";	-- 0x1D26
		when 007463 => D <= "00111010";	-- 0x1D27
		when 007464 => D <= "11001010";	-- 0x1D28
		when 007465 => D <= "00110011";	-- 0x1D29
		when 007466 => D <= "00111101";	-- 0x1D2A
		when 007467 => D <= "11011101";	-- 0x1D2B
		when 007468 => D <= "00100011";	-- 0x1D2C
		when 007469 => D <= "11011101";	-- 0x1D2D
		when 007470 => D <= "01111110";	-- 0x1D2E
		when 007471 => D <= "00000000";	-- 0x1D2F
		when 007472 => D <= "11000011";	-- 0x1D30
		when 007473 => D <= "00100010";	-- 0x1D31
		when 007474 => D <= "00111101";	-- 0x1D32
		when 007475 => D <= "11011101";	-- 0x1D33
		when 007476 => D <= "01111110";	-- 0x1D34
		when 007477 => D <= "00000000";	-- 0x1D35
		when 007478 => D <= "11111110";	-- 0x1D36
		when 007479 => D <= "00111010";	-- 0x1D37
		when 007480 => D <= "11000010";	-- 0x1D38
		when 007481 => D <= "10001001";	-- 0x1D39
		when 007482 => D <= "00111101";	-- 0x1D3A
		when 007483 => D <= "11011101";	-- 0x1D3B
		when 007484 => D <= "00100011";	-- 0x1D3C
		when 007485 => D <= "11011101";	-- 0x1D3D
		when 007486 => D <= "00100010";	-- 0x1D3E
		when 007487 => D <= "00001111";	-- 0x1D3F
		when 007488 => D <= "10000000";	-- 0x1D40
		when 007489 => D <= "11011101";	-- 0x1D41
		when 007490 => D <= "00101010";	-- 0x1D42
		when 007491 => D <= "00001101";	-- 0x1D43
		when 007492 => D <= "10000000";	-- 0x1D44
		when 007493 => D <= "11001101";	-- 0x1D45
		when 007494 => D <= "00100010";	-- 0x1D46
		when 007495 => D <= "00111100";	-- 0x1D47
		when 007496 => D <= "11011010";	-- 0x1D48
		when 007497 => D <= "01101110";	-- 0x1D49
		when 007498 => D <= "00111111";	-- 0x1D4A
		when 007499 => D <= "11011101";	-- 0x1D4B
		when 007500 => D <= "00100010";	-- 0x1D4C
		when 007501 => D <= "00001101";	-- 0x1D4D
		when 007502 => D <= "10000000";	-- 0x1D4E
		when 007503 => D <= "00100010";	-- 0x1D4F
		when 007504 => D <= "00010010";	-- 0x1D50
		when 007505 => D <= "10000000";	-- 0x1D51
		when 007506 => D <= "11011101";	-- 0x1D52
		when 007507 => D <= "00101010";	-- 0x1D53
		when 007508 => D <= "00001111";	-- 0x1D54
		when 007509 => D <= "10000000";	-- 0x1D55
		when 007510 => D <= "11011101";	-- 0x1D56
		when 007511 => D <= "01111110";	-- 0x1D57
		when 007512 => D <= "00000000";	-- 0x1D58
		when 007513 => D <= "11001101";	-- 0x1D59
		when 007514 => D <= "10111100";	-- 0x1D5A
		when 007515 => D <= "00101010";	-- 0x1D5B
		when 007516 => D <= "11011010";	-- 0x1D5C
		when 007517 => D <= "01101110";	-- 0x1D5D
		when 007518 => D <= "00111111";	-- 0x1D5E
		when 007519 => D <= "00111110";	-- 0x1D5F
		when 007520 => D <= "00000001";	-- 0x1D60
		when 007521 => D <= "11001101";	-- 0x1D61
		when 007522 => D <= "01110010";	-- 0x1D62
		when 007523 => D <= "00101011";	-- 0x1D63
		when 007524 => D <= "11010010";	-- 0x1D64
		when 007525 => D <= "01101110";	-- 0x1D65
		when 007526 => D <= "00111111";	-- 0x1D66
		when 007527 => D <= "11011101";	-- 0x1D67
		when 007528 => D <= "00100010";	-- 0x1D68
		when 007529 => D <= "00001111";	-- 0x1D69
		when 007530 => D <= "10000000";	-- 0x1D6A
		when 007531 => D <= "11111110";	-- 0x1D6B
		when 007532 => D <= "00000010";	-- 0x1D6C
		when 007533 => D <= "11000010";	-- 0x1D6D
		when 007534 => D <= "01110011";	-- 0x1D6E
		when 007535 => D <= "00111101";	-- 0x1D6F
		when 007536 => D <= "11000011";	-- 0x1D70
		when 007537 => D <= "01101110";	-- 0x1D71
		when 007538 => D <= "00111111";	-- 0x1D72
		when 007539 => D <= "00101010";	-- 0x1D73
		when 007540 => D <= "00010010";	-- 0x1D74
		when 007541 => D <= "10000000";	-- 0x1D75
		when 007542 => D <= "11111101";	-- 0x1D76
		when 007543 => D <= "01110101";	-- 0x1D77
		when 007544 => D <= "00000000";	-- 0x1D78
		when 007545 => D <= "11111101";	-- 0x1D79
		when 007546 => D <= "01110100";	-- 0x1D7A
		when 007547 => D <= "00000001";	-- 0x1D7B
		when 007548 => D <= "11011101";	-- 0x1D7C
		when 007549 => D <= "00101010";	-- 0x1D7D
		when 007550 => D <= "00001111";	-- 0x1D7E
		when 007551 => D <= "10000000";	-- 0x1D7F
		when 007552 => D <= "11001101";	-- 0x1D80
		when 007553 => D <= "11001100";	-- 0x1D81
		when 007554 => D <= "00100111";	-- 0x1D82
		when 007555 => D <= "11011101";	-- 0x1D83
		when 007556 => D <= "01111110";	-- 0x1D84
		when 007557 => D <= "00000000";	-- 0x1D85
		when 007558 => D <= "11000011";	-- 0x1D86
		when 007559 => D <= "00110110";	-- 0x1D87
		when 007560 => D <= "00111101";	-- 0x1D88
		when 007561 => D <= "11011101";	-- 0x1D89
		when 007562 => D <= "00101010";	-- 0x1D8A
		when 007563 => D <= "00001111";	-- 0x1D8B
		when 007564 => D <= "10000000";	-- 0x1D8C
		when 007565 => D <= "11011101";	-- 0x1D8D
		when 007566 => D <= "01111110";	-- 0x1D8E
		when 007567 => D <= "00000000";	-- 0x1D8F
		when 007568 => D <= "11011101";	-- 0x1D90
		when 007569 => D <= "00100011";	-- 0x1D91
		when 007570 => D <= "10110111";	-- 0x1D92
		when 007571 => D <= "11000010";	-- 0x1D93
		when 007572 => D <= "10001101";	-- 0x1D94
		when 007573 => D <= "00111101";	-- 0x1D95
		when 007574 => D <= "11011101";	-- 0x1D96
		when 007575 => D <= "11001011";	-- 0x1D97
		when 007576 => D <= "00000000";	-- 0x1D98
		when 007577 => D <= "01111110";	-- 0x1D99
		when 007578 => D <= "11000010";	-- 0x1D9A
		when 007579 => D <= "10010001";	-- 0x1D9B
		when 007580 => D <= "00111111";	-- 0x1D9C
		when 007581 => D <= "11001101";	-- 0x1D9D
		when 007582 => D <= "00111011";	-- 0x1D9E
		when 007583 => D <= "00111100";	-- 0x1D9F
		when 007584 => D <= "11001101";	-- 0x1DA0
		when 007585 => D <= "11001100";	-- 0x1DA1
		when 007586 => D <= "00100111";	-- 0x1DA2
		when 007587 => D <= "11011101";	-- 0x1DA3
		when 007588 => D <= "01111110";	-- 0x1DA4
		when 007589 => D <= "00000000";	-- 0x1DA5
		when 007590 => D <= "10110111";	-- 0x1DA6
		when 007591 => D <= "11000010";	-- 0x1DA7
		when 007592 => D <= "11111110";	-- 0x1DA8
		when 007593 => D <= "00111100";	-- 0x1DA9
		when 007594 => D <= "11011101";	-- 0x1DAA
		when 007595 => D <= "00100011";	-- 0x1DAB
		when 007596 => D <= "00111010";	-- 0x1DAC
		when 007597 => D <= "00000010";	-- 0x1DAD
		when 007598 => D <= "10000000";	-- 0x1DAE
		when 007599 => D <= "10110111";	-- 0x1DAF
		when 007600 => D <= "11000010";	-- 0x1DB0
		when 007601 => D <= "11111110";	-- 0x1DB1
		when 007602 => D <= "00111100";	-- 0x1DB2
		when 007603 => D <= "11011101";	-- 0x1DB3
		when 007604 => D <= "11100001";	-- 0x1DB4
		when 007605 => D <= "11110001";	-- 0x1DB5
		when 007606 => D <= "00110010";	-- 0x1DB6
		when 007607 => D <= "00010001";	-- 0x1DB7
		when 007608 => D <= "10000000";	-- 0x1DB8
		when 007609 => D <= "10110111";	-- 0x1DB9
		when 007610 => D <= "11001010";	-- 0x1DBA
		when 007611 => D <= "11010000";	-- 0x1DBB
		when 007612 => D <= "00111101";	-- 0x1DBC
		when 007613 => D <= "11111101";	-- 0x1DBD
		when 007614 => D <= "11100001";	-- 0x1DBE
		when 007615 => D <= "11100001";	-- 0x1DBF
		when 007616 => D <= "11111101";	-- 0x1DC0
		when 007617 => D <= "01110101";	-- 0x1DC1
		when 007618 => D <= "00000000";	-- 0x1DC2
		when 007619 => D <= "11111101";	-- 0x1DC3
		when 007620 => D <= "01110100";	-- 0x1DC4
		when 007621 => D <= "00000001";	-- 0x1DC5
		when 007622 => D <= "00111010";	-- 0x1DC6
		when 007623 => D <= "00010001";	-- 0x1DC7
		when 007624 => D <= "10000000";	-- 0x1DC8
		when 007625 => D <= "00111101";	-- 0x1DC9
		when 007626 => D <= "00110010";	-- 0x1DCA
		when 007627 => D <= "00010001";	-- 0x1DCB
		when 007628 => D <= "10000000";	-- 0x1DCC
		when 007629 => D <= "11000011";	-- 0x1DCD
		when 007630 => D <= "10111001";	-- 0x1DCE
		when 007631 => D <= "00111101";	-- 0x1DCF
		when 007632 => D <= "11000001";	-- 0x1DD0
		when 007633 => D <= "01111001";	-- 0x1DD1
		when 007634 => D <= "00110010";	-- 0x1DD2
		when 007635 => D <= "00000011";	-- 0x1DD3
		when 007636 => D <= "10000000";	-- 0x1DD4
		when 007637 => D <= "01111000";	-- 0x1DD5
		when 007638 => D <= "00110010";	-- 0x1DD6
		when 007639 => D <= "00000010";	-- 0x1DD7
		when 007640 => D <= "10000000";	-- 0x1DD8
		when 007641 => D <= "11000011";	-- 0x1DD9
		when 007642 => D <= "11011111";	-- 0x1DDA
		when 007643 => D <= "00111101";	-- 0x1DDB
		when 007644 => D <= "11000011";	-- 0x1DDC
		when 007645 => D <= "01101110";	-- 0x1DDD
		when 007646 => D <= "00111111";	-- 0x1DDE
		when 007647 => D <= "11000011";	-- 0x1DDF
		when 007648 => D <= "00000110";	-- 0x1DE0
		when 007649 => D <= "00111110";	-- 0x1DE1
		when 007650 => D <= "11111101";	-- 0x1DE2
		when 007651 => D <= "00100001";	-- 0x1DE3
		when 007652 => D <= "10000111";	-- 0x1DE4
		when 007653 => D <= "00110001";	-- 0x1DE5
		when 007654 => D <= "11001101";	-- 0x1DE6
		when 007655 => D <= "00110101";	-- 0x1DE7
		when 007656 => D <= "00101010";	-- 0x1DE8
		when 007657 => D <= "11011010";	-- 0x1DE9
		when 007658 => D <= "00000011";	-- 0x1DEA
		when 007659 => D <= "00111110";	-- 0x1DEB
		when 007660 => D <= "00010001";	-- 0x1DEC
		when 007661 => D <= "10000001";	-- 0x1DED
		when 007662 => D <= "00000000";	-- 0x1DEE
		when 007663 => D <= "10101111";	-- 0x1DEF
		when 007664 => D <= "11101101";	-- 0x1DF0
		when 007665 => D <= "01010010";	-- 0x1DF1
		when 007666 => D <= "00101001";	-- 0x1DF2
		when 007667 => D <= "00010001";	-- 0x1DF3
		when 007668 => D <= "00101011";	-- 0x1DF4
		when 007669 => D <= "00110001";	-- 0x1DF5
		when 007670 => D <= "00011001";	-- 0x1DF6
		when 007671 => D <= "01011110";	-- 0x1DF7
		when 007672 => D <= "00100011";	-- 0x1DF8
		when 007673 => D <= "01010110";	-- 0x1DF9
		when 007674 => D <= "11101011";	-- 0x1DFA
		when 007675 => D <= "00010001";	-- 0x1DFB
		when 007676 => D <= "00000000";	-- 0x1DFC
		when 007677 => D <= "00111110";	-- 0x1DFD
		when 007678 => D <= "11010101";	-- 0x1DFE
		when 007679 => D <= "11101001";	-- 0x1DFF
		when 007680 => D <= "11000011";	-- 0x1E00
		when 007681 => D <= "00000110";	-- 0x1E01
		when 007682 => D <= "00111110";	-- 0x1E02
		when 007683 => D <= "11000011";	-- 0x1E03
		when 007684 => D <= "01101110";	-- 0x1E04
		when 007685 => D <= "00111111";	-- 0x1E05
		when 007686 => D <= "11001001";	-- 0x1E06
		when 007687 => D <= "10101111";	-- 0x1E07
		when 007688 => D <= "00110010";	-- 0x1E08
		when 007689 => D <= "01001111";	-- 0x1E09
		when 007690 => D <= "10000011";	-- 0x1E0A
		when 007691 => D <= "00100001";	-- 0x1E0B
		when 007692 => D <= "01001111";	-- 0x1E0C
		when 007693 => D <= "10000011";	-- 0x1E0D
		when 007694 => D <= "00100010";	-- 0x1E0E
		when 007695 => D <= "01001001";	-- 0x1E0F
		when 007696 => D <= "10000011";	-- 0x1E10
		when 007697 => D <= "00100001";	-- 0x1E11
		when 007698 => D <= "00000000";	-- 0x1E12
		when 007699 => D <= "00000000";	-- 0x1E13
		when 007700 => D <= "00100010";	-- 0x1E14
		when 007701 => D <= "01000111";	-- 0x1E15
		when 007702 => D <= "10000011";	-- 0x1E16
		when 007703 => D <= "00100001";	-- 0x1E17
		when 007704 => D <= "00000000";	-- 0x1E18
		when 007705 => D <= "10000110";	-- 0x1E19
		when 007706 => D <= "00100010";	-- 0x1E1A
		when 007707 => D <= "01000001";	-- 0x1E1B
		when 007708 => D <= "10000011";	-- 0x1E1C
		when 007709 => D <= "00100010";	-- 0x1E1D
		when 007710 => D <= "01000011";	-- 0x1E1E
		when 007711 => D <= "10000011";	-- 0x1E1F
		when 007712 => D <= "00100001";	-- 0x1E20
		when 007713 => D <= "11111111";	-- 0x1E21
		when 007714 => D <= "10001111";	-- 0x1E22
		when 007715 => D <= "00100010";	-- 0x1E23
		when 007716 => D <= "01000101";	-- 0x1E24
		when 007717 => D <= "10000011";	-- 0x1E25
		when 007718 => D <= "00110110";	-- 0x1E26
		when 007719 => D <= "00000000";	-- 0x1E27
		when 007720 => D <= "00100001";	-- 0x1E28
		when 007721 => D <= "00110100";	-- 0x1E29
		when 007722 => D <= "00111110";	-- 0x1E2A
		when 007723 => D <= "00010001";	-- 0x1E2B
		when 007724 => D <= "01001011";	-- 0x1E2C
		when 007725 => D <= "10000011";	-- 0x1E2D
		when 007726 => D <= "00000001";	-- 0x1E2E
		when 007727 => D <= "00000100";	-- 0x1E2F
		when 007728 => D <= "00000000";	-- 0x1E30
		when 007729 => D <= "11101101";	-- 0x1E31
		when 007730 => D <= "10110000";	-- 0x1E32
		when 007731 => D <= "11001001";	-- 0x1E33
		when 007732 => D <= "01010101";	-- 0x1E34
		when 007733 => D <= "10101010";	-- 0x1E35
		when 007734 => D <= "00000001";	-- 0x1E36
		when 007735 => D <= "10000000";	-- 0x1E37
		when 007736 => D <= "00100001";	-- 0x1E38
		when 007737 => D <= "11111111";	-- 0x1E39
		when 007738 => D <= "10001111";	-- 0x1E3A
		when 007739 => D <= "00100010";	-- 0x1E3B
		when 007740 => D <= "00000000";	-- 0x1E3C
		when 007741 => D <= "10000000";	-- 0x1E3D
		when 007742 => D <= "10101111";	-- 0x1E3E
		when 007743 => D <= "00110010";	-- 0x1E3F
		when 007744 => D <= "00101010";	-- 0x1E40
		when 007745 => D <= "10000000";	-- 0x1E41
		when 007746 => D <= "00110010";	-- 0x1E42
		when 007747 => D <= "01000111";	-- 0x1E43
		when 007748 => D <= "10000000";	-- 0x1E44
		when 007749 => D <= "00110010";	-- 0x1E45
		when 007750 => D <= "00000010";	-- 0x1E46
		when 007751 => D <= "10000000";	-- 0x1E47
		when 007752 => D <= "00110010";	-- 0x1E48
		when 007753 => D <= "00000011";	-- 0x1E49
		when 007754 => D <= "10000000";	-- 0x1E4A
		when 007755 => D <= "00110010";	-- 0x1E4B
		when 007756 => D <= "00010110";	-- 0x1E4C
		when 007757 => D <= "10000000";	-- 0x1E4D
		when 007758 => D <= "00110010";	-- 0x1E4E
		when 007759 => D <= "00101001";	-- 0x1E4F
		when 007760 => D <= "10000000";	-- 0x1E50
		when 007761 => D <= "00110010";	-- 0x1E51
		when 007762 => D <= "00000100";	-- 0x1E52
		when 007763 => D <= "10000000";	-- 0x1E53
		when 007764 => D <= "00110010";	-- 0x1E54
		when 007765 => D <= "00100101";	-- 0x1E55
		when 007766 => D <= "10000000";	-- 0x1E56
		when 007767 => D <= "00111110";	-- 0x1E57
		when 007768 => D <= "00000001";	-- 0x1E58
		when 007769 => D <= "00110010";	-- 0x1E59
		when 007770 => D <= "00110110";	-- 0x1E5A
		when 007771 => D <= "10000000";	-- 0x1E5B
		when 007772 => D <= "00110010";	-- 0x1E5C
		when 007773 => D <= "01000011";	-- 0x1E5D
		when 007774 => D <= "10000000";	-- 0x1E5E
		when 007775 => D <= "00110010";	-- 0x1E5F
		when 007776 => D <= "01000100";	-- 0x1E60
		when 007777 => D <= "10000000";	-- 0x1E61
		when 007778 => D <= "00110010";	-- 0x1E62
		when 007779 => D <= "00100111";	-- 0x1E63
		when 007780 => D <= "10000000";	-- 0x1E64
		when 007781 => D <= "00110010";	-- 0x1E65
		when 007782 => D <= "00101000";	-- 0x1E66
		when 007783 => D <= "10000000";	-- 0x1E67
		when 007784 => D <= "00100001";	-- 0x1E68
		when 007785 => D <= "00110100";	-- 0x1E69
		when 007786 => D <= "00111110";	-- 0x1E6A
		when 007787 => D <= "00010001";	-- 0x1E6B
		when 007788 => D <= "01001011";	-- 0x1E6C
		when 007789 => D <= "10000011";	-- 0x1E6D
		when 007790 => D <= "00000110";	-- 0x1E6E
		when 007791 => D <= "00000100";	-- 0x1E6F
		when 007792 => D <= "11100101";	-- 0x1E70
		when 007793 => D <= "00100001";	-- 0x1E71
		when 007794 => D <= "10000111";	-- 0x1E72
		when 007795 => D <= "00111110";	-- 0x1E73
		when 007796 => D <= "11100011";	-- 0x1E74
		when 007797 => D <= "00011010";	-- 0x1E75
		when 007798 => D <= "10111110";	-- 0x1E76
		when 007799 => D <= "11001010";	-- 0x1E77
		when 007800 => D <= "01111100";	-- 0x1E78
		when 007801 => D <= "00111110";	-- 0x1E79
		when 007802 => D <= "00110111";	-- 0x1E7A
		when 007803 => D <= "11001001";	-- 0x1E7B
		when 007804 => D <= "00100011";	-- 0x1E7C
		when 007805 => D <= "00010011";	-- 0x1E7D
		when 007806 => D <= "00000101";	-- 0x1E7E
		when 007807 => D <= "11000010";	-- 0x1E7F
		when 007808 => D <= "10000100";	-- 0x1E80
		when 007809 => D <= "00111110";	-- 0x1E81
		when 007810 => D <= "10101111";	-- 0x1E82
		when 007811 => D <= "11001001";	-- 0x1E83
		when 007812 => D <= "11000011";	-- 0x1E84
		when 007813 => D <= "01110101";	-- 0x1E85
		when 007814 => D <= "00111110";	-- 0x1E86
		when 007815 => D <= "11010010";	-- 0x1E87
		when 007816 => D <= "10001101";	-- 0x1E88
		when 007817 => D <= "00111110";	-- 0x1E89
		when 007818 => D <= "11001101";	-- 0x1E8A
		when 007819 => D <= "00000111";	-- 0x1E8B
		when 007820 => D <= "00111110";	-- 0x1E8C
		when 007821 => D <= "10101111";	-- 0x1E8D
		when 007822 => D <= "00110010";	-- 0x1E8E
		when 007823 => D <= "00101010";	-- 0x1E8F
		when 007824 => D <= "10000000";	-- 0x1E90
		when 007825 => D <= "00110010";	-- 0x1E91
		when 007826 => D <= "00101011";	-- 0x1E92
		when 007827 => D <= "10000000";	-- 0x1E93
		when 007828 => D <= "00111110";	-- 0x1E94
		when 007829 => D <= "00000111";	-- 0x1E95
		when 007830 => D <= "11001101";	-- 0x1E96
		when 007831 => D <= "11110011";	-- 0x1E97
		when 007832 => D <= "00100000";	-- 0x1E98
		when 007833 => D <= "10101111";	-- 0x1E99
		when 007834 => D <= "11001101";	-- 0x1E9A
		when 007835 => D <= "11110011";	-- 0x1E9B
		when 007836 => D <= "00100000";	-- 0x1E9C
		when 007837 => D <= "00111110";	-- 0x1E9D
		when 007838 => D <= "00000010";	-- 0x1E9E
		when 007839 => D <= "11001101";	-- 0x1E9F
		when 007840 => D <= "11110011";	-- 0x1EA0
		when 007841 => D <= "00100000";	-- 0x1EA1
		when 007842 => D <= "11001101";	-- 0x1EA2
		when 007843 => D <= "00010001";	-- 0x1EA3
		when 007844 => D <= "00100001";	-- 0x1EA4
		when 007845 => D <= "00100001";	-- 0x1EA5
		when 007846 => D <= "00000000";	-- 0x1EA6
		when 007847 => D <= "00000000";	-- 0x1EA7
		when 007848 => D <= "00100010";	-- 0x1EA8
		when 007849 => D <= "11011010";	-- 0x1EA9
		when 007850 => D <= "10000010";	-- 0x1EAA
		when 007851 => D <= "11001101";	-- 0x1EAB
		when 007852 => D <= "10111101";	-- 0x1EAC
		when 007853 => D <= "00100000";	-- 0x1EAD
		when 007854 => D <= "11001101";	-- 0x1EAE
		when 007855 => D <= "11100100";	-- 0x1EAF
		when 007856 => D <= "00100000";	-- 0x1EB0
		when 007857 => D <= "11001001";	-- 0x1EB1
		when 007858 => D <= "01111110";	-- 0x1EB2
		when 007859 => D <= "10110111";	-- 0x1EB3
		when 007860 => D <= "11001000";	-- 0x1EB4
		when 007861 => D <= "01001111";	-- 0x1EB5
		when 007862 => D <= "11001101";	-- 0x1EB6
		when 007863 => D <= "10110111";	-- 0x1EB7
		when 007864 => D <= "00110000";	-- 0x1EB8
		when 007865 => D <= "00100011";	-- 0x1EB9
		when 007866 => D <= "00011000";	-- 0x1EBA
		when 007867 => D <= "11110110";	-- 0x1EBB
		when 007868 => D <= "01000111";	-- 0x1EBC
		when 007869 => D <= "01001111";	-- 0x1EBD
		when 007870 => D <= "01010011";	-- 0x1EBE
		when 007871 => D <= "01001001";	-- 0x1EBF
		when 007872 => D <= "00100000";	-- 0x1EC0
		when 007873 => D <= "00101101";	-- 0x1EC1
		when 007874 => D <= "00100000";	-- 0x1EC2
		when 007875 => D <= "01000111";	-- 0x1EC3
		when 007876 => D <= "01110010";	-- 0x1EC4
		when 007877 => D <= "01100001";	-- 0x1EC5
		when 007878 => D <= "01110000";	-- 0x1EC6
		when 007879 => D <= "01101000";	-- 0x1EC7
		when 007880 => D <= "01101001";	-- 0x1EC8
		when 007881 => D <= "01110011";	-- 0x1EC9
		when 007882 => D <= "01100011";	-- 0x1ECA
		when 007883 => D <= "01101000";	-- 0x1ECB
		when 007884 => D <= "00100000";	-- 0x1ECC
		when 007885 => D <= "01101111";	-- 0x1ECD
		when 007886 => D <= "01110010";	-- 0x1ECE
		when 007887 => D <= "01101001";	-- 0x1ECF
		when 007888 => D <= "01100101";	-- 0x1ED0
		when 007889 => D <= "01101110";	-- 0x1ED1
		when 007890 => D <= "01110100";	-- 0x1ED2
		when 007891 => D <= "01101001";	-- 0x1ED3
		when 007892 => D <= "01100101";	-- 0x1ED4
		when 007893 => D <= "01110010";	-- 0x1ED5
		when 007894 => D <= "01110100";	-- 0x1ED6
		when 007895 => D <= "01100101";	-- 0x1ED7
		when 007896 => D <= "00100000";	-- 0x1ED8
		when 007897 => D <= "01010011";	-- 0x1ED9
		when 007898 => D <= "01110000";	-- 0x1EDA
		when 007899 => D <= "01110010";	-- 0x1EDB
		when 007900 => D <= "01100001";	-- 0x1EDC
		when 007901 => D <= "01100011";	-- 0x1EDD
		when 007902 => D <= "01101000";	-- 0x1EDE
		when 007903 => D <= "01100101";	-- 0x1EDF
		when 007904 => D <= "00100000";	-- 0x1EE0
		when 007905 => D <= "01001001";	-- 0x1EE1
		when 007906 => D <= "00100000";	-- 0x1EE2
		when 007907 => D <= "00001101";	-- 0x1EE3
		when 007908 => D <= "00001010";	-- 0x1EE4
		when 007909 => D <= "00101000";	-- 0x1EE5
		when 007910 => D <= "01000011";	-- 0x1EE6
		when 007911 => D <= "00101001";	-- 0x1EE7
		when 007912 => D <= "00100000";	-- 0x1EE8
		when 007913 => D <= "01001101";	-- 0x1EE9
		when 007914 => D <= "01110101";	-- 0x1EEA
		when 007915 => D <= "01100101";	-- 0x1EEB
		when 007916 => D <= "01101110";	-- 0x1EEC
		when 007917 => D <= "01100011";	-- 0x1EED
		when 007918 => D <= "01101000";	-- 0x1EEE
		when 007919 => D <= "01100101";	-- 0x1EEF
		when 007920 => D <= "01101110";	-- 0x1EF0
		when 007921 => D <= "00100000";	-- 0x1EF1
		when 007922 => D <= "00110001";	-- 0x1EF2
		when 007923 => D <= "00111001";	-- 0x1EF3
		when 007924 => D <= "00111000";	-- 0x1EF4
		when 007925 => D <= "00110100";	-- 0x1EF5
		when 007926 => D <= "00100000";	-- 0x1EF6
		when 007927 => D <= "01010010";	-- 0x1EF7
		when 007928 => D <= "01101111";	-- 0x1EF8
		when 007929 => D <= "01101100";	-- 0x1EF9
		when 007930 => D <= "01100110";	-- 0x1EFA
		when 007931 => D <= "00101101";	-- 0x1EFB
		when 007932 => D <= "01000100";	-- 0x1EFC
		when 007933 => D <= "01101001";	-- 0x1EFD
		when 007934 => D <= "01100101";	-- 0x1EFE
		when 007935 => D <= "01110100";	-- 0x1EFF
		when 007936 => D <= "01100101";	-- 0x1F00
		when 007937 => D <= "01110010";	-- 0x1F01
		when 007938 => D <= "00100000";	-- 0x1F02
		when 007939 => D <= "01001011";	-- 0x1F03
		when 007940 => D <= "01101100";	-- 0x1F04
		when 007941 => D <= "01100101";	-- 0x1F05
		when 007942 => D <= "01101001";	-- 0x1F06
		when 007943 => D <= "01101110";	-- 0x1F07
		when 007944 => D <= "00100000";	-- 0x1F08
		when 007945 => D <= "01010110";	-- 0x1F09
		when 007946 => D <= "01100101";	-- 0x1F0A
		when 007947 => D <= "01110010";	-- 0x1F0B
		when 007948 => D <= "01110011";	-- 0x1F0C
		when 007949 => D <= "00100000";	-- 0x1F0D
		when 007950 => D <= "00110001";	-- 0x1F0E
		when 007951 => D <= "00101110";	-- 0x1F0F
		when 007952 => D <= "00110001";	-- 0x1F10
		when 007953 => D <= "00100000";	-- 0x1F11
		when 007954 => D <= "00001101";	-- 0x1F12
		when 007955 => D <= "00001010";	-- 0x1F13
		when 007956 => D <= "00100010";	-- 0x1F14
		when 007957 => D <= "01000101";	-- 0x1F15
		when 007958 => D <= "01101001";	-- 0x1F16
		when 007959 => D <= "01101110";	-- 0x1F17
		when 007960 => D <= "00100000";	-- 0x1F18
		when 007961 => D <= "01001000";	-- 0x1F19
		when 007962 => D <= "01100001";	-- 0x1F1A
		when 007963 => D <= "01110101";	-- 0x1F1B
		when 007964 => D <= "01100011";	-- 0x1F1C
		when 007965 => D <= "01101000";	-- 0x1F1D
		when 007966 => D <= "00100000";	-- 0x1F1E
		when 007967 => D <= "01110110";	-- 0x1F1F
		when 007968 => D <= "01101111";	-- 0x1F20
		when 007969 => D <= "01101110";	-- 0x1F21
		when 007970 => D <= "00100000";	-- 0x1F22
		when 007971 => D <= "01001100";	-- 0x1F23
		when 007972 => D <= "01001111";	-- 0x1F24
		when 007973 => D <= "01000111";	-- 0x1F25
		when 007974 => D <= "01001111";	-- 0x1F26
		when 007975 => D <= "00100000";	-- 0x1F27
		when 007976 => D <= "00101110";	-- 0x1F28
		when 007977 => D <= "00101110";	-- 0x1F29
		when 007978 => D <= "00101110";	-- 0x1F2A
		when 007979 => D <= "00100010";	-- 0x1F2B
		when 007980 => D <= "00001101";	-- 0x1F2C
		when 007981 => D <= "00001010";	-- 0x1F2D
		when 007982 => D <= "00000000";	-- 0x1F2E
		when 007983 => D <= "00001101";	-- 0x1F2F
		when 007984 => D <= "00001010";	-- 0x1F30
		when 007985 => D <= "01000101";	-- 0x1F31
		when 007986 => D <= "01101110";	-- 0x1F32
		when 007987 => D <= "01100100";	-- 0x1F33
		when 007988 => D <= "01100101";	-- 0x1F34
		when 007989 => D <= "00101110";	-- 0x1F35
		when 007990 => D <= "00001101";	-- 0x1F36
		when 007991 => D <= "00001010";	-- 0x1F37
		when 007992 => D <= "00000000";	-- 0x1F38
		when 007993 => D <= "00001101";	-- 0x1F39
		when 007994 => D <= "00001010";	-- 0x1F3A
		when 007995 => D <= "01000110";	-- 0x1F3B
		when 007996 => D <= "01100101";	-- 0x1F3C
		when 007997 => D <= "01101000";	-- 0x1F3D
		when 007998 => D <= "01101100";	-- 0x1F3E
		when 007999 => D <= "01100101";	-- 0x1F3F
		when 008000 => D <= "01110010";	-- 0x1F40
		when 008001 => D <= "00101110";	-- 0x1F41
		when 008002 => D <= "00001101";	-- 0x1F42
		when 008003 => D <= "00001010";	-- 0x1F43
		when 008004 => D <= "00000000";	-- 0x1F44
		when 008005 => D <= "00001101";	-- 0x1F45
		when 008006 => D <= "00001010";	-- 0x1F46
		when 008007 => D <= "01010011";	-- 0x1F47
		when 008008 => D <= "01110000";	-- 0x1F48
		when 008009 => D <= "01100101";	-- 0x1F49
		when 008010 => D <= "01101001";	-- 0x1F4A
		when 008011 => D <= "01100011";	-- 0x1F4B
		when 008012 => D <= "01101000";	-- 0x1F4C
		when 008013 => D <= "01100101";	-- 0x1F4D
		when 008014 => D <= "01110010";	-- 0x1F4E
		when 008015 => D <= "01110000";	-- 0x1F4F
		when 008016 => D <= "01101100";	-- 0x1F50
		when 008017 => D <= "01100001";	-- 0x1F51
		when 008018 => D <= "01110100";	-- 0x1F52
		when 008019 => D <= "01111010";	-- 0x1F53
		when 008020 => D <= "00100000";	-- 0x1F54
		when 008021 => D <= "00111111";	-- 0x1F55
		when 008022 => D <= "00101110";	-- 0x1F56
		when 008023 => D <= "00001101";	-- 0x1F57
		when 008024 => D <= "00001010";	-- 0x1F58
		when 008025 => D <= "00000000";	-- 0x1F59
		when 008026 => D <= "00001101";	-- 0x1F5A
		when 008027 => D <= "00001010";	-- 0x1F5B
		when 008028 => D <= "01000101";	-- 0x1F5C
		when 008029 => D <= "01101110";	-- 0x1F5D
		when 008030 => D <= "01100100";	-- 0x1F5E
		when 008031 => D <= "01101100";	-- 0x1F5F
		when 008032 => D <= "01101111";	-- 0x1F60
		when 008033 => D <= "01110011";	-- 0x1F61
		when 008034 => D <= "01110011";	-- 0x1F62
		when 008035 => D <= "01100011";	-- 0x1F63
		when 008036 => D <= "01101000";	-- 0x1F64
		when 008037 => D <= "01101100";	-- 0x1F65
		when 008038 => D <= "01100101";	-- 0x1F66
		when 008039 => D <= "01101001";	-- 0x1F67
		when 008040 => D <= "01100110";	-- 0x1F68
		when 008041 => D <= "01100101";	-- 0x1F69
		when 008042 => D <= "00101110";	-- 0x1F6A
		when 008043 => D <= "00001101";	-- 0x1F6B
		when 008044 => D <= "00001010";	-- 0x1F6C
		when 008045 => D <= "00000000";	-- 0x1F6D
		when 008046 => D <= "11101101";	-- 0x1F6E
		when 008047 => D <= "01111011";	-- 0x1F6F
		when 008048 => D <= "00000000";	-- 0x1F70
		when 008049 => D <= "10000000";	-- 0x1F71
		when 008050 => D <= "11001101";	-- 0x1F72
		when 008051 => D <= "11101111";	-- 0x1F73
		when 008052 => D <= "00110000";	-- 0x1F74
		when 008053 => D <= "00001110";	-- 0x1F75
		when 008054 => D <= "00111111";	-- 0x1F76
		when 008055 => D <= "11001101";	-- 0x1F77
		when 008056 => D <= "10110111";	-- 0x1F78
		when 008057 => D <= "00110000";	-- 0x1F79
		when 008058 => D <= "11011101";	-- 0x1F7A
		when 008059 => D <= "11100101";	-- 0x1F7B
		when 008060 => D <= "11100001";	-- 0x1F7C
		when 008061 => D <= "11001101";	-- 0x1F7D
		when 008062 => D <= "10110010";	-- 0x1F7E
		when 008063 => D <= "00111110";	-- 0x1F7F
		when 008064 => D <= "00100001";	-- 0x1F80
		when 008065 => D <= "00111001";	-- 0x1F81
		when 008066 => D <= "00111111";	-- 0x1F82
		when 008067 => D <= "00011000";	-- 0x1F83
		when 008068 => D <= "00100111";	-- 0x1F84
		when 008069 => D <= "11101101";	-- 0x1F85
		when 008070 => D <= "01111011";	-- 0x1F86
		when 008071 => D <= "00000000";	-- 0x1F87
		when 008072 => D <= "10000000";	-- 0x1F88
		when 008073 => D <= "00100001";	-- 0x1F89
		when 008074 => D <= "01000101";	-- 0x1F8A
		when 008075 => D <= "00111111";	-- 0x1F8B
		when 008076 => D <= "11001101";	-- 0x1F8C
		when 008077 => D <= "10110010";	-- 0x1F8D
		when 008078 => D <= "00111110";	-- 0x1F8E
		when 008079 => D <= "00011000";	-- 0x1F8F
		when 008080 => D <= "00011011";	-- 0x1F90
		when 008081 => D <= "11101101";	-- 0x1F91
		when 008082 => D <= "01111011";	-- 0x1F92
		when 008083 => D <= "00000000";	-- 0x1F93
		when 008084 => D <= "10000000";	-- 0x1F94
		when 008085 => D <= "00100001";	-- 0x1F95
		when 008086 => D <= "01011010";	-- 0x1F96
		when 008087 => D <= "00111111";	-- 0x1F97
		when 008088 => D <= "00011000";	-- 0x1F98
		when 008089 => D <= "00010010";	-- 0x1F99
		when 008090 => D <= "11101101";	-- 0x1F9A
		when 008091 => D <= "01111011";	-- 0x1F9B
		when 008092 => D <= "00000000";	-- 0x1F9C
		when 008093 => D <= "10000000";	-- 0x1F9D
		when 008094 => D <= "00100001";	-- 0x1F9E
		when 008095 => D <= "00101111";	-- 0x1F9F
		when 008096 => D <= "00111111";	-- 0x1FA0
		when 008097 => D <= "00011000";	-- 0x1FA1
		when 008098 => D <= "00001001";	-- 0x1FA2
		when 008099 => D <= "00110001";	-- 0x1FA3
		when 008100 => D <= "11111111";	-- 0x1FA4
		when 008101 => D <= "10001111";	-- 0x1FA5
		when 008102 => D <= "11001101";	-- 0x1FA6
		when 008103 => D <= "00111000";	-- 0x1FA7
		when 008104 => D <= "00111110";	-- 0x1FA8
		when 008105 => D <= "00100001";	-- 0x1FA9
		when 008106 => D <= "10111100";	-- 0x1FAA
		when 008107 => D <= "00111110";	-- 0x1FAB
		when 008108 => D <= "10101111";	-- 0x1FAC
		when 008109 => D <= "00110010";	-- 0x1FAD
		when 008110 => D <= "00000100";	-- 0x1FAE
		when 008111 => D <= "10000000";	-- 0x1FAF
		when 008112 => D <= "11001101";	-- 0x1FB0
		when 008113 => D <= "10110010";	-- 0x1FB1
		when 008114 => D <= "00111110";	-- 0x1FB2
		when 008115 => D <= "11100101";	-- 0x1FB3
		when 008116 => D <= "00100001";	-- 0x1FB4
		when 008117 => D <= "11011100";	-- 0x1FB5
		when 008118 => D <= "00111111";	-- 0x1FB6
		when 008119 => D <= "11100011";	-- 0x1FB7
		when 008120 => D <= "10101111";	-- 0x1FB8
		when 008121 => D <= "00110010";	-- 0x1FB9
		when 008122 => D <= "00000010";	-- 0x1FBA
		when 008123 => D <= "10000000";	-- 0x1FBB
		when 008124 => D <= "11001101";	-- 0x1FBC
		when 008125 => D <= "11111001";	-- 0x1FBD
		when 008126 => D <= "00110000";	-- 0x1FBE
		when 008127 => D <= "11100101";	-- 0x1FBF
		when 008128 => D <= "11011101";	-- 0x1FC0
		when 008129 => D <= "11100001";	-- 0x1FC1
		when 008130 => D <= "11001101";	-- 0x1FC2
		when 008131 => D <= "11001100";	-- 0x1FC3
		when 008132 => D <= "00100111";	-- 0x1FC4
		when 008133 => D <= "11011101";	-- 0x1FC5
		when 008134 => D <= "01111110";	-- 0x1FC6
		when 008135 => D <= "00000000";	-- 0x1FC7
		when 008136 => D <= "10110111";	-- 0x1FC8
		when 008137 => D <= "11001010";	-- 0x1FC9
		when 008138 => D <= "11011001";	-- 0x1FCA
		when 008139 => D <= "00111111";	-- 0x1FCB
		when 008140 => D <= "11001101";	-- 0x1FCC
		when 008141 => D <= "00111011";	-- 0x1FCD
		when 008142 => D <= "00111100";	-- 0x1FCE
		when 008143 => D <= "11001101";	-- 0x1FCF
		when 008144 => D <= "11001100";	-- 0x1FD0
		when 008145 => D <= "00100111";	-- 0x1FD1
		when 008146 => D <= "11011101";	-- 0x1FD2
		when 008147 => D <= "01111110";	-- 0x1FD3
		when 008148 => D <= "00000000";	-- 0x1FD4
		when 008149 => D <= "10110111";	-- 0x1FD5
		when 008150 => D <= "11000010";	-- 0x1FD6
		when 008151 => D <= "11001100";	-- 0x1FD7
		when 008152 => D <= "00111111";	-- 0x1FD8
		when 008153 => D <= "11000011";	-- 0x1FD9
		when 008154 => D <= "10111000";	-- 0x1FDA
		when 008155 => D <= "00111111";	-- 0x1FDB
		when 008156 => D <= "01110110";	-- 0x1FDC
		when 008157 => D <= "00000000";	-- 0x1FDD
		when 008158 => D <= "00000000";	-- 0x1FDE
		when 008159 => D <= "00000000";	-- 0x1FDF
		when 008160 => D <= "00000000";	-- 0x1FE0
		when 008161 => D <= "00000000";	-- 0x1FE1
		when 008162 => D <= "00000000";	-- 0x1FE2
		when 008163 => D <= "00000000";	-- 0x1FE3
		when 008164 => D <= "00000000";	-- 0x1FE4
		when 008165 => D <= "00000000";	-- 0x1FE5
		when 008166 => D <= "00000000";	-- 0x1FE6
		when 008167 => D <= "00000000";	-- 0x1FE7
		when 008168 => D <= "00000000";	-- 0x1FE8
		when 008169 => D <= "00000000";	-- 0x1FE9
		when 008170 => D <= "00000000";	-- 0x1FEA
		when 008171 => D <= "00000000";	-- 0x1FEB
		when 008172 => D <= "00000000";	-- 0x1FEC
		when 008173 => D <= "00000000";	-- 0x1FED
		when 008174 => D <= "00000000";	-- 0x1FEE
		when 008175 => D <= "00000000";	-- 0x1FEF
		when 008176 => D <= "00000000";	-- 0x1FF0
		when 008177 => D <= "00000000";	-- 0x1FF1
		when 008178 => D <= "00000000";	-- 0x1FF2
		when 008179 => D <= "00000000";	-- 0x1FF3
		when 008180 => D <= "00000000";	-- 0x1FF4
		when 008181 => D <= "00000000";	-- 0x1FF5
		when 008182 => D <= "00000000";	-- 0x1FF6
		when 008183 => D <= "00000000";	-- 0x1FF7
		when 008184 => D <= "00000000";	-- 0x1FF8
		when 008185 => D <= "00000000";	-- 0x1FF9
		when 008186 => D <= "00000000";	-- 0x1FFA
		when 008187 => D <= "00000000";	-- 0x1FFB
		when 008188 => D <= "00000000";	-- 0x1FFC
		when 008189 => D <= "00000000";	-- 0x1FFD
		when 008190 => D <= "00000000";	-- 0x1FFE
		when 008191 => D <= "00000000";	-- 0x1FFF
		when others => D <= "--------";
		end case;
	end process;
end;
