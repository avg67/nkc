--
--Written by GowinSynthesis
--Tool Version "V1.9.10 (64-bit)"
--Thu Oct  3 21:53:41 2024

--Source file index table:
--file0 "\C:/working/_Tang_nano/_cores/ps2_fifo/fifo_sc_hs.vhdl/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\C:/working/_Tang_nano/_cores/ps2_fifo/fifo_sc_hs.vhdl/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
LCnl6cPN9tX1PSxXqcUtDWQP9o4QnCCrvIvoxy6Wctia39fbP+rA09jm/WSjA5NnvshfVCboNpsm
7BY/C0XvnfUL99esGDezEzbjF9Q6/7zMWp6S6c2swDzJAZ38dmqd/6ATmrJPu+R/ad7hzhqmLHOu
jMrAE1btWHWfsnUhxUJ+h2Tf76izgGlRJPGV0BsJvq9GuLia56Xx3JAG2tFvvIe1IzeYYGLhXnBM
L6yGQTmf+e+LABIXWjDehEiFoAHUBOfb8Pcwr92L2oEu5Twju1r0bof3tgTy37ovwihc4wKbdItA
UZNtQkWD81lI3wTBsLIZVqC8SnCo4qUSaJIULw==

`protect encoding=(enctype="base64", line_length=76, bytes=53840)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
Xh54CiFlL35B2KEIQjiaFky/Ww5qOyy8NuFkx8Nd2TZYRm5f+v8KH2qe9xFDmCvKvFRY6tx7GuTc
NEHkq/T972PMV11kfZhKt4NMdBmECv5B+KC2orGpWjAiLW1XOM8fGQJOkaFf2q5oTkF4lhyVcYK0
FR3n3zPDH0uvyFw+oxKLTDiwmimnzY8b6D9hN/kg0++eHa91PGWtUcgJmYKnM0BBA1v9Lz46lpB2
sFc0Ed5dS3gz164lebK+PKSe1ymMSk+sJn0j3m1nD3lFfzWfPKuWPKIG/flGSp+sDsLIBHbQHzg6
lNuK7mUBRvT5LacEc7uLoV8MRjPltUPigty1HSR2hrpA2Xa6yGAKK71U8zkbbnsxIA+lO8ik+4rq
JvOiQODL59SQGBuGZXLw5KeDbwwUnJXHSkVRgDdtLCVninh/NxQkVouASbIZq2Lr0tzc2w1ptH8R
V9ljPRMC572y9NgUGXyerFENv4dZiqe2rt5ApiWQ18MOxambUQWP42EM3/PwQaScsiiCDHAALbu1
Bqgb9Qv8mBaLM8fLBVcrGaNJ/1/xK6hIJNFi4CxhEotc/mcbpc3qk9bxaB+ejC69TxsZ85xIH+Sg
lsJO6s0ge9DkSOZC+6vd2HVzsPyjtd5RZvodRulhwBG/ryaFDChwE+fGtEYSkJIVFZAbF6UkwheQ
XGKie85kzERedeUMmQunuHvMffNHG4lvu5uJq1GC2g1M7Iqzi7j7kBvDUS+QX/uo0KaSwiH+XJEQ
GqmGTxA9ahSzX4KHRKU9LyQVpdjiQsRD8ZWpE/nRcpqv1frMrxRkerEt6GVrSjtV/fBfxn531bNe
9+pfogrJtTrzPTzlW2eYweA7mlsHOaOHSFQqzc47c8tOVhUp/oowwt002nnTQCu2Ui2TUj5UB8fi
4Mz8p3PbpVzeygxO4s6uPIDtIZbDIrNmHNXMJGR9s+eJdZfwEzYoT08UYJFab02O0L0Gx/EHjr3V
EG0IrcOBV60L5ffxQiwcmHQYbgJINDt9iqKNGHwylArMW3m5g9HK0DD/M4gd3F5FKBBtu39GbZJz
SS9Ml52YXgxDe5FLEgtYzQcr8lcpfbCZEIKPzO7cyBg+HFI9MtX5Bxai3EllmfZ3vJTZ6kTyZ1n8
czV4T2QKALrzdhCSJr3z+ix9WfQ88guxMUKsXD84W4v5VteHeKwUOso/klwDnIYC7Vn1kiN/sSJz
z//x3g5GuPWQ4cgWt4ou5B/2Tb9OVXySS8gl+bbadRVV5gysKEBEGTsOTXr4mOrjezPyI68w0eYb
JyKhYtzZgzo7PaZn49WIhpgVnKyz3BHoYY7aENhBg5I+jjAj3CzCq3SeLsu/EVRd8UeHVyML/Wjv
zdHe0Q/Nh6U1cVjQNUeZqUG0/mRLq5xTeh0RXDzccyqers3uXKbGb/1sZz1kPFlttfc0yi90J1MX
MMx2wuzDUWhDvxwqVZXOXCtMb46g+52CB5CQjZU0/TOMsF3NpCNvHAZ1q6NJUOZOVdMiNWmZpZl/
wgIdGcoS0uAH4vpgVTqSsXnHqgvPPCHI4WtlhwIPms4Sb7HE1NuWYum1qxE71xhKaHw/7Xnd38kz
DNp8zqKR2BJviHuIZLLOMrKfc5eVZf0LotndUyKT/jF2aa7kuYHJR07E8PzL+cUqbchAQfNwzf5J
Z722iYq/i77J12a2YWMu1wsvH57SALVPB1jzp4RUUelheAT3GpYnCqr7kcRBpjiutx3SG7RPHUP0
4CjMsW7fQ51sGrDy7wWmNrYEKENRwVnW1LqXlYClThONGWJQdGDdKsVleZ0RMOPHydd0xlmPT85B
7Lc9ba9pCkfPgY6Hdlzl0SQMHTIzLGwHNDA8uwNePbeR6dly/50jONcd+x8BStNl61XBW7KwGUtJ
BUTL3UOqjeuJV3itCSjPnsqoaFYu7ooZgeVu+7eoQDdlmIAJ5j6Rt03nnnBxxU6tO2Pp2fChzgJR
wxa6R41Ymku61Pzz92Av/n68PKr8iSafdk5TTGGDlKP9DK7gFbCeJZBudt4WeP1i+PXj/urp/fcN
XfoPXcNezOd4npEEx1jtaHMeJn/HHtW6QcNdK65It/lkRLHriyxCWHme1WtuHlwKTPMSWSDV8zHD
dF0c12UvdES+lqYEdssPTZZCftPNJn0cyQl85EZXZsI7MkfFhZ0AlTuVi8D2GeWS4kzLyZtY4yKQ
7QyY9fYCo9xHtqP3DDqIFaOOgRcHxwQzeYCBjaZgj5rdAtcJhibLnLHpH/FAwqMCYbISp6sihRDG
5CMMAT+h5E2bhakmyyMiNQk47COZgcdo0c6637nJktKzukznWi7cs+bIEOJypeLUivBqjPEJtq4i
5UYPkokI7NRMdEKGetAy90tRdQKIaYC+qO2BkSSJ5zBOk9RNW2e4lO3tTIkWw1AulSAA5KCP39o9
ASha9LAsGqA/4ikxzi+u/T0EK8epP+3i7BUkNf4FRNxDXcAVsN9Vp69mF5odTDT0tXhNGwrZEJml
SkbTiyfQNaQ4MZpPyijAsubalA5yraHnIf9bXsi53WjlqNAb5t44unNZTfYCZcr5h24bSyBG/BQk
B5LOm/uDE1o36u7k87Jubfaaq63iA8Zf3cb4FQ6KsTe9+Zb2dgDMGmDKzAojLXZYE0pUDMH9EVFc
Y/7qIv+Um5oDmf9Zdr+WMnlxxim2IWVAqDirQB+mBcKk8Fa6Yd/NsdbA8i5pKjaFe5gq4ILQOyjz
8meZRFeelJG8IgGPqcEgOo76bAsYP1bDLSUrsLwljju2gqsW33ppzUkdbJ48Fi6pVkBpUwoO1Dst
lOG3qfhfqUZy3dZO98KfPWiLxR4PB7W2p1qdDKZ1oR92L+e49WEHFqaYZu0IhceXSWJDKo52pJnO
DwQAeapI8B5dPEPioQHpUsJbIqiDADezUnlsJ6EZNPf11dN1qxf6ZvU95oPzKgkpY4hecSYy0EO8
U6SOG+AqhzhKqbUZLxzYibjdbVqkkY2O9nRJ8C7gHCH4ON+PvnmRRz8wZ/K4wdi9203rjJE7SZqt
SxXmGRNCYHtHquT8sLaTusTn9whmLsFJ5VY9lC0LRJOGwLIjwfyRdkSRPZgZhNGLsjTdwzlM1utr
U77C0/e4FaAHjUiFik/gdBy0Z/PNOwljUjDUYOmjUtDz8kyWfK4bTDH1l4clgHB2yEPzK4J7qV39
K2UUWr0SAH5QFVxRcMYMf+WUd7HBfZJV+9CpJmTlGBY0R86vWzCrzz0dnVcDDECweaAfqzfr3gVA
FgQUR+0c0nPYGNE1niA70evhrzR1XGogRhy0dnIjNwQhGP6D5hjPR+E7C9BVFAmQa6O2ptZA7oLI
nnUId32c7q26XSm/z5byX/yjAiLQ+YI5E37K3ccct7s4uvCliKwgcJx5Ib3px/oTTo3vUBoWrRNR
tnjLV6i6tEHUvV8kH+Z0ZdRMi/pUZOAG/QO/k5v4BN/fBuelVENea2BYjhK1jW/04BxV6/WEEWOX
EBpjJdWjABAGCqQRT8qmT4MPfyKxK1Rvff5HGiZtS9TYdN2R5iDivNADMzQYBHhw3XX1rtzOQ/fZ
YreFOuITheT2sLiZWrQG35J/Q0OM0LhL3OG2CJj6VTGYEYflvRZuOyokzJsHXAQZaMv/Zh7PaFkE
8RJLo4qGvHQFT+jlE5P71KvygMdsnpVB5JIqTVIOHNApoYZ4SrZr/NjMr2FQJ5ksSibubJ6sw/ED
lgrtwiHeabA5NYgmnhJNUPCBPOHnDr9Q/Cs5UHFQNp9wYBY4AF5o5fteigAaPiaZrr38M9E4CYEk
ViwkDvptHSVsaQO1rTETk44T+cd7cVRpji9ebpx9jYjMuT7FqOifD2RU0yznW35RodsJ67Ha20xm
RV1pj2WY6i8GX5pR7UJp0KuXKk82mCzUydAJ/EUiR6OB2vKw1v3xfD9XMzhpnuRfEFi/d2k011Fy
no5s/0o3GeW/FQb0Uzw6V/66w2w0Zsh2aNu0llXnhIuSUXfSwDpfICI5a82ZRS/o9/9KbGp71zw2
1v++kbaLHBP/IMT6HzXPpKY+1qDPJLBsgKJtgYFNWK98DfOOdWhmtAJAI5BQ6wp9CcFJyM51zaik
JANyxvWehNghCg5B1X1bGolCtrqDB0X5/pcP+nFXTB9FxLj/0XY8lRaL3BSx12yMXYPFP+fmLrqC
WaPAuvDSHRhS46fPKIEJAskyrqbPYZ0kZiSIaaYdVYiAcrVJKLvhaJhEs0kjFm0EujtJUVjVXUA9
5E/IaDuYa1W4uxrwZ/9D43Dg6SdGEL8t9PZHqhdrev7o3U2tz1mEVWNEhsS0ekuLZgI76jHc6Uz1
nzrGTEUfoN1l1P9uVg3m++eJ3NAls+oKfBl2PCL7gQeGJD+JSbVTCX488O8egIbrOtGwsxccf7Sf
gdQWiAornP8MQkP+q/p+6ODJr/oCMu2fW9K5Z+ea52flqOKmiWYr2cgyPQLRuzYDmrfSDE6gwAho
3XKhtzjjPOWSIDdWjTKmkhB0gWYHnvSneGkiPe4WefTCjIB+EuEhW4LAuyhnGQyn61tZ90ntONyU
SnNsIecS8gwno8B0iJKtiEc1EmZGRqrZ97ahhiHC8H9HUHneKYx1+h/UFCjqc647skah1YJyeced
uzu1kZUknvE6IXs7OGpP2sVtKqp4TFSAggx8cae4HnAOGIqnTkNbu0t5YtRnm2Fo5arUdurwT55+
c6hYvCMCwLUCi/okNESJFMfDhyC5LtFExKy5VfJhtFc1WYxWGxbX4fFs9lsXU44CH4JMchQCeHv2
kRnBRjPGqLLCUliWSaNdO2ppUSqb9tk5pTuzlY+XNcyrVOYBUOQGEdaxESYtFFhdBzov+93o04NO
dfauZrMR6yA4b4qbi2qOTL8rn4bDvrfrBYioBnlK8XTpT8ZzLDnv8pxew6zQyV+B3E640jfk283P
PrEkrG5rGO4zpQ++CC8WDs0LYdHGJZp6/xQCjNLdoqFj61mDjcTm9djSwmKNPwfW0FLY1ApGs0rI
keCHZAtWc5XGCZoh4l1BNjFgofqssrakrkYcFYX0ZPPa3NMA+8OsgJ1d+d4GktZImv1YL3Sr/rm9
xDtzsnv0ZUGPyny14MSAcl1bc/VW2GTSQdzZn0c9odlfU4Caq4i9tEB6xBoXDVVRRF9gNvWJdOGV
g9azP4qx2ToNgALTv8Y7ZemHCcr3zkpsHaCeg3ye9R2wiV17vz1f2j78ZrT2wUr/+8F3Zbe7LmsD
PPcP/93nAi8Eo22LyCvvwOe1/rj+gEjbSI0p4s6VFpziIgzBE0PAmpEOn+g1o6AcpzPBjzssnJrU
qMYSgAP6pdXaILa0QCc68LnsMvMTq7ubGEuHOWGqowJdfFVmnAH1zQ5JH1RKAst1uFlE4eDdQOkM
WdeDNa9Rlmr3vdN/q0tEpf27zpWsygvJSkoYg0OuK/o56lC7NVz0wiCuqd04apW1kWFoxvKfADbQ
nhWGdh1C1DSCxdD4OzTOR1ioyIy+MDBvbHthc4N54Ao3DkjwxBhm+ZsOwit7CHH0duJWw9/i24qP
iB5HwuxDELU5ytfRpamu+K8WqMc1g+9crR+JbPbNpWwgZvjCrGh08fRQ587ZJjspZ01kK9dPfSqi
hu2L59btXVpOQJqMaTxxw0TMkd9xTult99MZVVEmK85aRjwZFmGIz3veEBzaRP2Aeo/w+8l/ZAen
0cWF+QC8OtvYuNGSTb/nOaQkr3G1rP3vm64rLHXI/maK94lF4RwxKpng5JZU5DvTwj+azyqvfttH
MzpvpcjK78lRjbDw6mjjzuB867iOHIub0TsR9XgFf5gPmIC93ayj/gFi7ucX6Ks41BjYI2rpBTWW
LsSLr/phvElFc85ZH8liSzwQXvtkuf0TnYLhOW6Zoh797gB8uBVdDlsTwuv7SBN8mvJFkLUYWkBQ
3vEf9OZMjUMKd7oM43QPGHgzIjQN4ezlRcGOCu2MLfkyGSRCNGjWV1i66IbtGUEkdgjf2mSYwNaf
F741ezuhKosUQ0wi6UzCfUC/6v7NLcDlJZSl4KwHqy9Bpg4iqlQo12egqmuCyILjR64myc8FjHGj
4FuMXepSadzRxaO7oOSI3tojPUGsQsAdOZhOgTy2QHhANAPTkATkwk4BLAq0wF7VpeawCL7GD88i
ZFY6yQlKQAoWzYxYmxBoRaXmE4GKwoeCg2OfRQu/Hunt6IDqV7DFTFxzuxa2Ffmi6aNn8RczvF2I
4bbOBRJmW3fKyp6FpUtfbBh+i2aGX0K/XKMXKnQPtTnK3u6sqDD91QdGm8BoxWXNUOyBiC+R6Ag8
5/g2y6dczmmiSDk7+irlPyoSY6D6Ig4ZllIzseIC+UvTQM2fwsYaHNi6W19LFunEzu2oGIeeiz//
WLSfV6R0V66g17HguapAGUm34dIo+Bw+/iU8LnUBQakK/uxG88GFVQZ2xqXdwV+sv71rNQOyRcru
0mRyP8zXU03jWarPkWSlmdhhUwKsJFqYAwcCQKPeUlk/G6h0TJ84WpM9SM9Z2alqFlBom5E9PRw2
h0wcSro1GveEYu03sbjC3c5XpRtgZxI04y1rupJm+GQzOI6myANSaUfNZs66hl3UXg+YWN3bGi2/
UptjJVAQoH07hp2tz0MZD1/Z0CwlSnRfTIhTieH6T+IpGz1hlfxWxU/lmUFKb/cS6MUE/Q5iLuV1
vhqul9VjZ0hTYvPCwEa4AimVel9H2D16Sq3ujqqCZw0hq9YnbzrvoPO8eQyLzdUVtKE8D/mKI5L9
xJ0//LrnqmuN86mVHKKZ2Vz0QLK5I2c8G8UsVHp90YCVxvbQ9Wa4Er6WKxy9FomUjmhTKviXrVd3
WKNFMi5Tsl6p6dvWjJfbMsKX5M/eBtrQQ/Dv6d7S66L2vauovV92RbHSZ+6UvjV/UN23zCN1yNba
h7x/k5XGt/HkwVcKvaS8Q6MpUGGC8qAMSzPP7wnCYyWOGdB60jAIy2WCXz0VGt+JkBfqhweQpjx8
qgO+5T6mBkNzv378MiNf+fvTQ73Mg++VIQhC5j8vVqECIDW8vc++bZ1psijOYbWshywy8LOrSimx
ZLN9lFr4IXPS12NEoTjIH5QQhQK8bG8DFtyuDZnQDG92SiOpaiTpNNW+uaZP1zU1VguT0O/2MOYD
rgTjw/S4EmJvcpST5VWfdXfknxUVfw6dxoMIcKXrEIGo6mFvq5zbGsZ6e/5ylDq+cgfn3Cc+/2HE
4ETNFA2OTBRm6nnQRLr/wMmDbJCzUh6ZvpvamBuIPnzaXKGi9AV3nkP8LHv1/yzOkdfTRch3joFZ
IToTshZCu1NtbOrWqxlYP50cbBgjFk66NTTzwd5Tg4XzAXl07ezR9N8kQKt52mcTbedSdgbTUXc3
iDiixbQ53yVUUyK0R06Yx1Z+ktOLBKUnv8yHii+cMivkVZEC0qLUF1907SGJBwDD9hO/wKS6SHUy
dMZpvV4yvx/6GjO8lu8mWRRsZRuLidHS5sKJlhEUxxx5E5z5TNg8WFl5dM9t7n701zWysTHMeugZ
fYvUvGAtcm2gdngtZuBI1wWvH07E7JzFR1hNNTjD7giUCz3JqcfpgTBnIvmn6AruRL6lEzs2moHB
wCoym5PNnVCfEEd2W9Tq29Qj1EuZCPp6j9hQH8/MjqxNfx9vXJCROMubV5Acgg/XtqvmBqNnN76g
q+GcqNjy1+JgWhQOgf9gyU1/EkZjhTXdkWUrgWe5BdC7yduHQpb/xM0NcmIuLu59pWb/l2mXgHp7
v4B6BT0OFSaH+qfYx1PNCwm99x2k62Nyr9rrWVJVSR+lS5YzTIfHffdo2n0ykTtAC3Icps7B8Inr
a1vUd0Oh/4FDeQbmTTMRpxj9CkG/0zfy8Hl0yzo5jjGdSAAmVw9a5ja6r+vVBOr4hWuIGa9jM9PJ
3ZUUvIOydt5pp/PhOT5DRoXVcB3278KPGHfxsaUkr4ChCPib+AQhe7F2Zq32n0aW79BrL6M4f6pB
+7vvuWPzw3mFicBCZ6DR19ev8fiuqCSQmNTBpAjPRcCA1c+Y5Z45JfYfI8N0trxW7vs+tvj2nGoy
JNWoHnUn/+yuNZfAU/D1rQ0crT6Yuv+z7s+7Oudoe2OQL/pHzZinPUDOyuB7+3EiAjhWhLoPs4YB
pncmaUSpZnyWos9ajKLt4/I8IU/ECGFH1//024p8q+/aVh+HqWZJPwL0nuJnfpzfrZK2g4Q9lsB5
TYAB9uXGka/dNvq8THvpv5tyMuYY2hKwf+J8hH1Ke/KOji75oO7P+Ye7NKSZNaoONSeRFMxv4cz1
lxgkgVkbw8YCD9VGBp4dS1EFYtf7Cb9vRYnn4bM+KTVPkvVDLglNfDIoLStKdd2hGhptdBPJbS0h
8jjp2rsW80WEGYyrQHThrgiOLAEvuegeFlGsi6rPe5jsD1w+1fgRKRLxZ0HgQwVdymEBpG549OMY
0Z+WMfoFGhExYte1FDEIa7feZJdNjzFVSCzZeq1+uil7qx9bh2Eq26prKrMyJGQBtSAgQDG6nAfy
iFrk5C2Qv6X9xUQQlv6JvNQS0J8gfvIhGiFjO9GZwWaOUpV9Flp2tGARRBqOhtPWMEp5RtA+CmMl
N8SPKs3I8E19wfRYXOuHEwUkxZnhAXUTIW4Vc16DAkSL7+lT87fFcGsfBGkQxu8rO8jKub2VsP/I
sBnWxOc05JT6NFNhlePaDpXHwi8Mw6hC2k5qnmHEkvVYMCND36/YaIZQzqaTX8dnoiWVhf84RZjO
8p9k7gujTEPtLGrs0KLRjGBXY7dHxRSy5+qg6VPMQsYFl2m5KHzRrnFH7/wbDsdQK4OEn0PBWpsJ
o5qScB7BSkDAAM2DG12HKQ6qnaT4x3WNVFPMGLfG4ecCeKmEfRl98YMm8xxKrfT1q6Jae++ixTCs
9qnfwQhwbaXPJOMI/3Pa9KOK/bBpakZpEthtgOvm94VGpQdfdt53GjmstBEMChy7+sLsJq6LT4nM
R6pjQIxfjxQw9s4dJH5lINLzDz6ayZWVR8ur9Zmcb/PrGsNBbzTrspLvA9Qz9OWi38aFGRVgOChu
Og31lUIdz//11dpF0JeHKuwB02lny31BkunFADvB+ersM7ucTeu6jYOTffSmr9z9wGLVWzSkc+Bt
PhDrdDFZ3bi6x9AH5eP2fvw8f4rVrXLFXN7Nt2JfDZ188mUIMU0DGqNdhAhtlEAdZD1xwt8apkpZ
sbLKlAP5GQrz9rveMmKGtqsDKwTKrIda4mD3JqpGCCEQxTx++EcmQv8x/J+JqvgFox+UHAPmKVed
nCp94dt5VZcvuBG6mK/6ZaPvqJjafaIrfs2gRpvAkYAz9tc+QgBY4beePix7xW1D2tFCafsbCx4H
gMkKdeohT5xo3Aa2tGp0fkzUSC+N9zpDSFKWg3de1rXhOgNnH1Yl0ryU3lAZa/vBa7HsBDI57c+h
xhiZ4rXFMZB/b6VacvuEvLlE7VpDPLOFdHBk9/SQabVMv+tJ64HWhCXHUVLQfW3ymL+tae9lm/Qk
Bo5p3psVqLzoHSPePhb9OtTjWm8t2PL/Va6iJVsODZwYTPpDTHNQb2r3g47wmzM68yqJWu931Fhy
EPDA4BGEVk9pyRtpIKSKGbMVNzGGY/wX4XxEFD6xYPCyYIu9YU5Dkg/dIlwChLm3Q/2SQtKUwh1g
4Bd2mokGREvqOy+OK6R/ajANn6kimgNDqqcdLKJBLXKerq0vB6bfA12G9ExsEzyXndyAmnRn4DJt
vu9s09O96lWonuLUWqZK0k6XeacYY5y+UGbJCI1NmlFd7/fW1qYmX3dQ+otysbye4iAD7CwJm5cC
+bpY174XvHebIIQb0eUpIwRRSm/jbkBhyfIPoH16t1tl9imeLZh+xho468O5vG7eSmuG2CnTNC6E
CcXu3MDNSNaziaBi4PCMnUyrPGMWUvauVP3baEtXNICWz2NvsLcH6Q4i0dllgarDQ/hgQWEUDCu/
Cyuc1BwxubZQhNCae1jSzoB4mgVmXWoNu7wm6v0lfQyjcztzS5hBc8hUNadyfxG/qqKkDePCsICU
v3lg+W/EioJrSHo446mH/xXclJ/5lrsjK6L0QyaddiiD1QhBjxUgCMhkzE9BY63EgBOyJcLqwdl3
99HYmtZ35+jk0q6KgK7YcRDGMc4lEhGfmm20hPv3t7fRVn2INZ2MR9s03+hw/SRExfEbxHVh0/iD
27Kiuw6DN3u32pauadyirgzcqE6TlDkzj/HcHi1TKf++tndHEvN6EgUug02LVxI1e9tkWgh6rnM+
GB2LuCiW3k8m5AZnn31oPfXH6Kl9mVIC8QKLvMm/9rLJqszAGnNX26L17RAB23LzILMFjL+VO7Mf
FJPS8frbxC2tu/aIx04Nh9yc1c1/gr/t15rZ8ZzI7nyDW8zXhZ028MkIxCm3ndwpepL5knoOI+1B
26WRx5gBEF25JF5sCm7oqivxZA4mYjfWR1UIvlElyc8Zw+ok3Ke1uMcTnIH+aZqSh7cwNQ3xBn7p
XpaKqWz1ZjTnQ/FGxsvZqP6u/AViUyqv36hGR3f5gE6pxWOmHBGOs0vpxllXotZIr4/WUFO4yu1t
8nWI7KXx8imcgnlCN5yz2FnEfkrtk39h/yosNFYmDDIcKj3Bm833Xngf64/Xg25Ko5+X/7q8Jpc+
lKfV3Ozw/xlzrGjJNkYNPk4NYCbXb63WEohDXuuD/GtcMf6BTAIir30y0zsrgeCm32QvFqkjpYGY
jTL4xRLRWM8KcWS6PpPljPV8mdJUF+bHXPljbVPs1F2giIIx0tH/20FaimvLPHpw+bDQTU6qF8NA
JGMz1Mol565oSAsbu5FkpqEf2zkjsxLQqLBXROxMlotIbZ//7PvfDQ2xZ9BSLO87TZ7st0wpd/w3
+RVl0oApkGws1v4aM+43cXK9qx3Jgmsr3qyRWGOoYPbWEe5hPgyLF9qWDABXWOS8K5iEO+QmrcFn
8IzaBmb2UdcFbQNsROfa/4l0DSmB+lqaHRZUdb9wpFaolX2ftC0WbHZHywihPtLXV4n4mj6eGPbW
/ixLBwL0EuQeYvpIUcg4FSWlXancoPNPkJ5ycNXvwsNk6pi/7eUSHObB1YoS7xp0xdUZ1xWMa4E1
3zTiGfhJoAgKcjO+nRVhdzOuWFSBMFH8iiW++7W6mlBiMUcDu6pFDQL1FcXOnmz1ORt2e7nOPhiH
fZih31IZ+pOf4gnNwLlS9ZIq6NqspSe2FdBDZ+5axw6ZeLXO0AeZ0noZA5rgmDJpE95ySJb5ACFp
cvDAxNx7gXhmUlpAAYDf7fwmmjTkgK9hVuK3s0+F8YY0ywFt/3F0uaVOdbaD2L/vIgdpmv9BqazH
wTs3mc/C5xqzX5aDynUY8O2N0rP7YjMlO7yewPrY+JlY2EKy9TSCDRhRpmbxkMZy1GBkOGWUnt27
fWbBxwBNZmCh1VK87x9s0J3kieCcjPFbm5Cq3Vg8hSKNgF4EoGlto30uiCps6pk0Otw+3/LJDPUO
nrh6D0cwrxZqy/TOzeku3MVOWkSKqu2p6fVyBxVzZ7kUqwc2TP528tEBoPt2My1VXYXi8atXurSZ
JrTANp6JIYCIQd7zyiPbqx3BMUnzrXGG70OFUITkBRdgPQwTiA6qygRl/xyHc0iGjR719CEp01zw
6UWiNg8fOPSlsdlxmlrsfntWb3qmLKYj/6jrJO3p9YmFHI7OtTDkcrcr85q8M35pk9AL6UQIspJl
kThJG0h6pedl5lqWhNsQeK5ScuD4ioBLB2zVbK444UWReZQJgiTzQ+N6xykbWzVFjcjOXi6dngbY
0yBCH5UUQDInhKV+j+N1BywzCVl6Tc27f3zZQioi1xqtxg9DqV5LoCeMt9nbGGRXWXGZOglyDvWh
2J6V76txiOnUMO+RuhsO6RtALALiX7khWjM8PfeSNvMOS/V1u8GqxW/QTT/YMBwyD3+SFNf8wext
Y/ZxwQZnfWxxtdMDqzfpBtzo0mdwtviKki6DXJrlYPZpwn7sOxKXKEhwwv0bav1LU5o2s1ovq1s+
Kco1Nr6S4x7zy42WEprTUGV/LNb5hVsIeVJcdHhdM90KHRJbS1+t+8xe83U1u/PlMunJ5A8cWl48
g8MxUZH0K7C2/UvUSQ4mFvbYcylwadoouuLA4Z8xjmM5gBYKjby78dFTOHGNMIy6D9qLvrTWgQeR
OdgwCI+n+gr+gsI5qLzgC0cJRY1awwC7p0RZzSziC6yJWabCQHxCABgkgqkK5OK3akG82l9cT21b
ydaXNDvQkHHmbtvr4EK3ZEYtMZU5dJCwrYajPSLpKnhKH3bqdowvVZ0XSIXTNuYyKkWyb/iB2qCD
OAiKeEP3UtTMlhx57QyKMRYN6XD924bW/JwSGP5gGbvrq25joa6eCPfDEJm/hjvcdTSibqT1n3Gc
iSdBeg70mLC0q4+hT4J/LrH3KDfMn7wcO6cPC+3JpD44z30nYwJhaL5iMBj9x+yo/RJ+Rmy3I+V4
cQymK+ojF6k0HiZ7MoraYf7R9L/69kUpAr8j6/xi5xTbrhS/aWq7DAYAbaTX7F5ni296NzUWnSwh
hC6J81Hk73AcEim4GUs+TzgYRa2hclSxjvWWHeHEussPjOtjOw4wN4q95+Q/fBRE7pCy+poTcCK0
xvMejwEH/pa9KnfofvNdyvkYoUnOX20wTG409cYCHdRckYjGy4ZoZqLEwj+HozW9q+yb+8KINC3f
RQ75FCxys81+eZJ9MAbrtJ+feFWOwM7Q9ZSGpip/67o/i8uCwAEoCGRJp2XR+znXBYWqjJisM59V
uj1BXUdoDzRwSjCO3BXYbyWXCTB87mmrEDKhHmyldVcMaofP+8tAEPIn9ue0uxLj+5PqGTh+3ixh
jgnoxD4ftkTKkoNlu/TFXc3VqP3idv+REX78z9CKvsLCRhFaTNmbd38OzMyOIqhYeFIT1Re6R4ot
hwN1YgL9iuVDvWhCnSaBmp84mJ93l7ObRZzAKXI1fZOG+SoTHMxIxyI/2RSFwiKNDkQY9bJCrp+M
j2I/foJ/DmrUVKq3saxMyvYVI5RuYvaCUV5npoOK1MVWrfJsz8bMPST0YJlc7spDShrupPxPnTBV
JdSE9Kvxi4+7yVwWDLBxwGNd/oCrJ04Lu5UeI2/kCb3Q2NgR2tmNy+xI7ZiNt3fFA3I2zJ762sVl
0iYMSXM6TvEZsMZqkaQUd9wX02bWcBCtNBTdBdAavvGch4mq4nEHLq+EDzeOjjZP2zg6mcuQAGUr
RkBTuRnAlEHip0i09Rb4Y4+LF7nuRsoFlLF9fVoEzA1fxe9j+1AFcGIFA2CgyUZ2q9XV3/g3ncJB
7D1Qc7xDkUWH714u8G+he8y395yszq2tFfvSCnU/xhEglAjrh+Sl1ws0yO+U0sj36f7eR5XR6XHE
jJ+aYA8IB+CsCps77u00bfm66H4/Xi+QcxIIkkuKVir2Odw9hH8aBIyi38hIuy4ACb8EAgs5X+Ou
5J63n6xkWzdD1oIYymmqJyR7QMy9LkeQB6ZwB+GFFHI7lBIfaioVVoKym/ebQFDf0QHEDUi8Xct4
U2IAAico/j15ySEiZtBtM80tVKBZEspKf/17qAVpRr9MGc1OUyjfYahO/rLfUtFonhu2Mcw16CD8
zElAS3DO5ECzU1j3/qIWgsnA5M4FLHKsKbqAG1559aYpZZ8+9SG320dbqN1X9F+VDtnlWwemwj+v
GaHDCRuRwPbMm2lsT+98wFwO3HayTYrGq2VPtugiy24Dv/ZoJHqQu8Z3XuWDbI3RoGY+TTA1iVHY
GxGhNWcpigqVr+DfZBM/eRfvXcrep/irTqYbkCgp/zjlJbEdur92VIMktU68+NdQ2+lDbMvRuNI+
YGmcu2YN/9IRF+Vxwh0o7f6lKKA8FdRQ0l5l+B7xWP5hSPOyn6dKFCtUOAVNbWo8oNNJlItfN5tR
IucbJNlCIxucTLErjHHgrjN48/wNQv2Q+jG8PNYGvobVQ0G1wzhs7QYEnacDWddOytmK4p9K2LCS
cOCODLYaPyHBCsB1xIo3dQwwIFVSSlOFeCo1G66ArpyrzvgUUVkOR1YuHFVCDXnf/16YWvvTM1JF
hRiC6q2Yv/iNTqlNJNdh7t8shwKSYgy06X6JkESBRvP1v00dY9VZMzzgn8uV2CwCXBeB9Rl1MuXb
C/f7pSVSrGPHhrc5sPikutAYIJBwnSl6JAhIla4Q5HL2Je2P5+qFJ6C89Xey4A3AIh43zjz6cTZq
+8fvse6Aea7SWXZfk8/ay3u4kavx4y/DelhVoMQYYCSED7onlElZLQ7OYmDkxUyD/TZWVAwsdyjE
cmiLoBLwH8vRdYcpyGOFgAaHiYrXWoxdIpItxyfD6zdu7zjcZqxvbEZ8uuQLCj6G91rEMkPcqbHp
h+xeL/3L/ahEJLYgQeB2XSQKt1rroh35oy7mwScJNRnjSfTJMdS7ldj5CfLBV7oc0kVxCOm6HQOU
MOKew1wH5m4fpbLbngKPUxC2FaLPRb4uqRXTqSrgLSSkIsY1Q8hZgGALYAilqo3WBQ+4jtdju8dB
uNfKL0O+KZ7queh9LO1v2/Hnw3hUn8Q7o0kGbEXMCvDqVbgrzP98IEyKu0VTZOVP5f2vfzucIMuO
MoVcbA668MLWb2xJJntw+DpkoPZ5+1Z+mcUisAEl8CDxrdezsFJw8WV+A8t7x20bq6/9ch215uC3
RrnqN9TJfj14EDJOgUXS4TuAG32BpimbmmcmPgijGUsdfXbOlF94mj9Q5PSizeSF1L5enBv6L6nj
zuO6lEMe5z2Lqot1eij7RkB5uorQ4CjFWGFuoHZCvZhOKpCvDxHBFcfgVvAyOFzEBkZoVUNMVXzU
uD+4FeJnM5GdgLezYNZdsLK7IBsGfE1KKl7/0qiVKFOn1vOqpTQ8QLRcP7u/gYlui9M6eAQOq8LD
lZtG/UeDlS0IQ7kIFfDdfRGTYYItePG5Wjbupgzoo07uZn8SQ/rt2WdMrvp2QJL3vVxTRwxE58ir
5v3ObcKxsIeJxZ4Vj6B9xukX2FHeoesoP1OnolVwijMCtfpJGjpsMfRcGNN+LjaWqHEHHBb4N+8A
hibo683U6wKb7nPQDyMU2G5wPehU327YNvlhOj15vkLYydanbWllh3hSnLma2PRqNhDU3KyzOGY0
NxPo0FksfmSyIx3g1WOvTmcvyVwxcxgVL5kg6R4ig09BXVys2YgHtTxmL4vSE70mGCNOUqlhPnXo
/L5bCxgBSXvlbKK9IqR1j096zDb3fhHtrRvL7p0z3bFAML6UfRQHWNq7vRH9c/EGwUtvoiZ7XeYc
H1llTbpYasiJv6OiLPFi4PQxeP9WNhIO8KGJgdxk1vR6ALcHVRg8rscwMA+HxPXj9Im8OtQNMPt7
0aU2koQr3WWlrad7BRPl0KJTEpkfu1UF13WPdN0rP+rnbSLSi6fXg2P2XH+Kcw3LKU8iMTEFwsPL
UuekEW77JvsT4XxtNvEQDHeOGZvvpn00MHS4sF3UZ5BCv7XohO3UZFCgVOYvXozBoQtiH4DxixJG
m4bz8uzEFZt+33iGoNXemduCP+4tMzXPG7apmhhL6vzPv2m5IvMgcEGcYSZyCwc0ukXdkUl8nVM/
Jt9OCYGn5g03qfyXBcISClXReoByMYVGqvkJ1GIHlR4dfErSqf4iH4JoRpvxmfT/Zx7jz0PSxEyC
4JDFjqdG5O1pw9K3cmKwmMNKZQ5bQRvFhIXDxgl3alqfOzE36EHjwAkH2QGLGE+Z8hh7jLvgy9Yb
HH2cNZmZZQMPEAtjeek8wq/57du9n20/lw6aW64v3fYt7Qc0N6V5dJCdAJRfH4UIKZS2nROkgNU/
LKIghnBEgVJqZi7qhaobJ5uVE4VP20t12JZdj2UQAemYOho6vhRQeMU7zAltnTJoh2YzGD9pyQ8n
FhWxSQ7UsSGry9tdxEbt3oyVBjk+I4IUUEf+0Yxg3wqPHbIJWHHuKSrnQ6Z4LneLhAEVZl9J8vCc
cEthVQTt/b33Io8JnSol8u/Hi0I4PkfiyZ5qqY/k88Pe7rYXySoyQs8c3idl3MU2oMtuLi9c5k8/
LStbMUDZoaVCxE48CL+oRKTlBAob15YlC5+aCGzQiNToJ/Ww7e4r0JDTm7XCuqGQhpg/GqYXJodv
lIeoA7OBO9CNh7OrGFBbtsBInJ5B5JtqCoY5qLOBt5huSGp5IK29HXY7qv/qXmHdEompqyWDBZ/8
L3fIEgcXa8YSshirsCLZJQZxOxInE8TZH9TGFw/lfZ/mzRhankO0yKaPbu/Bu+N9xiIuNqbR6xzT
Dtkq/UaFj1dhZqWm/1oP381QV02aZEVA/TeBOhhhMS4VgXMNZiyre/Aw3tvo1BV+Wad8FksWTH8A
eg+6dL24UeNp6sUiNW/aJHO217oosL41YorSvWpE0YvpI/t7P4bjyR1JW5H10rOP5vH+1obrYm8p
ydnJUaiNO8UYL+4txHQRtlFotzp2vMpdx5751EqoVKy0bb0Bt5ZHgWzKC73eXRxwn3Xp030u5BK+
JZZuHaix8KjhvBQUV/kvQdvl/JudOe6tou1eu7fVF+9MhwIkgRuqtGTYpjNruOIQvCNK8BOWp9fD
v2QlAk/8fw6Fw2Qt8xL4RWO79/eC/OrN096lS57rom1x7TXDZw0husSjB0m7gdkvLy1si64tR4B/
WTd8UkJg+bvRFEoFYQgpqbwbXyuYNCOgSXRrorUz82GAVexBJHGPB2ubrm0tsQlT5niybABLutN6
sVupscDY2653z7rgefXPoL3/r3Qq4IqmqCMaKYAZdhA0kQHbs3C7AF7NZ+98+6fisQCv3kw4tEl1
YT+7OrNV88fHdmHE1+L4G32D72M6yVgr2qLYNMXOl+bFO8bPokI3RqwF49hT/W8rP2m9Pw2VweE7
8Qi9seV7vl6ZktXJP/oaxq8nAW+5ZJYCPFiZS0YEdLA/DwzIxcQngNn4UQ8OI9/WIQb3lgVMcJJo
L97p6YEgXsgpbd2iH4vO9FxHPkKH2q7iyWxK6pKc4hveOpNuj+dYas8F2LPW2xJausrvTFqej11h
4jl4VMXpM0xJcYzojzbgsANdRGNFcKHwx+fRxe7X/a/1JuvHRVljmF5KxuApJ3vdaUQKn2/Nh8G5
izLQ31e4rHWslcSIc56tV/72QstjPkf1Kn8LZSvf51SkZOdyPriMJVsEOjuY5wEEaCEoIRuwcWXZ
yqlg2HMjuFeGv5IzU8OBydmPdptC3D5rDY1v/bGzqYxmI39en552MvLs66zY94T3OldjOJHFsNNP
i9IGBkHsvZWQjn24lsKV0RFxMpmT42ErBkQ/zbKgFqm0dTwL/mQtKkiIFoE5lEMoECwfxucjU1D8
DAu1q99uKGHMtVTmBY7JWNL9u7WsM3k2evzMgUwp9rpkQoAM3PYHyPbEnclEAlJrjhF/sCZYyV+3
EMd+XJ57Jdm7YmCl+jJB3XfS2LSnuXT9ucC0n12pYxeyFo1MYk6PeBJ8tYp2LOdB6440uSxRelvQ
XPKMdJIqRiT4+6qJGBMk+72+oEu/S7Fr4aetN3wsZYzdbLtitoSSwWC9zIRuvyFOSk4QDNJUI/pA
pBfwH+ZPgrDeNqb5AfSeoDjqHF0XWRWrFbPdogKoAH+sgTWsOA63OM/bLNJn6TQ9lD4uU2ymDvqM
nEDrb7AYQ0h2qlNt6Zjo4FCGLPjSe/ibhyIAfqf5YsgLMZor6NaWFB3WKvatizni65H8ABDzeqfT
BAxY92eunBUIuQ1lbHjVu5TB0zSEKAUeneyZE8dJmuRe6V+7qXKIxruJ6iuPD2IYLC191BUM5jNh
uRDny5cElZfRM7bGvzlbdHhl1MgvDFC67ZVj1AHsCk0K+5Qq+v3r5I4Tx8/BZxm9N0h5sKdK/zqf
9oQZagO1IwINjuVr1nrRKc7hz2RU1ONgLqP6vvT+YbPw7lHdRFUMjbsjmpRC+l7qIFsVkhiPJnm8
42ZUFAyqmpzGcV/GUTNvLiZFZqUfbioi3Mq5ipSdDbouGM/Aa9Pn8b42OriSckMrBTPayL3B7l+6
+G8AHbMzl9k79PGxjszHKXQVuTYZhKvm1jE28RqG9EjKuf+I55ysfkbLddgjBZBmKxkpaiM6nat4
zEME/+G+2fPTgbYzElMuLhmTujsihTRoRYRZNi04mIvGJUo/ymTktlv7qP69bMsyxzitUQ5tFQzW
v/gIkP3AK9PACQXEXm+vm2EOWJARCkkLtC/DIDRI3WJv7xVZv6FnJa3MFKGMf8wkQAx8/o8LtxKq
DT6DGsO0DSXWlzyc701G2xDWw7QX3qriGS0x9OQXcbIX5MeTrzgBOvAYa+IqBmLhRPv0SYTk8Thd
GzQ+P5KRkPB/Jc+ErrYuGrxRLXDUnU5Txb6MuyaLR/G3GmRHKnQQeZNfRYtSTFntrUYmjOomN9BZ
XiSDihOXzOVcCAnyPhof/UIAPrHeC20iH9vWpnAd3cw2aTxIrFs/6YdNLpdzDH9poYkqUzScZavr
uFJy/M/kQAEImdsFWsCHuyADJXgX/53PrDzID4+BN9gsN/baAS9RQSkBCg66eBipG9hQM3XKZwgx
YpQfpGHlc5KUXvTXasYaEeM6nMRRZ0xa3zTx1wtPehJ0ZT7MYAgqLdg+DrTIPK8hM+bYSuirmgJU
EQ/Dz3BCROj6fZyJ/DT8MgmH2UAy+zqE3igK74hHwe6IV2qRBLxxKZ+IOwat3ggY2moQS+U3nICv
PcFBduJMejZRVRWV/L43GTHk271n4buyO6Uwv5ykqAZ7ulf9zUKGmWh8ZzUoX1MlDF48Q8dx6l2B
7aIzsLm/BH01ITBQX6LtGwacydCOfeTLn4O3I6J+8teFzMoYtbVsdzIS+4cG0wXGooIcB3cVVgUv
8I+sydSpd/rq7pz7fHiL4U/0aT1lKgf4N+79tpgU+tF9Bf2NWwwMDk0E2P+fHrVBx0mcFPPblP/S
fs1r+CB1zI6tbB8xtulkqiGIuPJytzMUzOE9SPb2e4DK5Z+u96pKKUsfvPcXI1Sxs4Yrf1klrk/1
GJVOla9Lu6yqg0nAC52a+WIltH0qt9KC31hYWy8dbSHzt4UsVRGNKLWOsmSkDllQa7zYMuKW6xSx
fpq+0WzW9XlA8fFPsb0DHuxBIyICShbeOBqORjesHYtUsQm0suWf0K/pmgYqBWd1+POI3Ojip7AN
OuqxEPqx3cp7q4r3BUM1qGBYKnF+zT9NBlSunrvWBqewvA2wxigY6G68mGoN7tqR1sR9pnRUw+za
SRVfhrfYc95eWFdOHgviarAcoKfGJexATIWPnoER7PVWdraHTX9xPh10jYRoW4eo3f+G1lm6LOOU
/rE8isd+ty1ibGa8O0ISDkx+YSuNJvBEWKqGZLnICKIHXZlT4Rh5EYe6bjNrVVAQ7RWYMGIG5yx/
AqNNX0VCXjtaglX67ZYbeMV4sXfRzxyLIEhpLRvdu58LOs0wi6jfiJAvQqA8fpBMGgplYXrt6Mpj
e9m8so6uyEU6UBX1rZQEIu5APYJhhHhOx0IxTeg0PENMrx0U9UrMHYQcwtMTjpZrua2UDjCxMDR1
vsj863XdyN0rc0dX7sCptA3r6OKS0/nMR8PyRdX7mQBPOH5A0O4m4CA361wZ2+mK1lbxw5ktATtN
ZTYwXhrEwQBx8vZblYTu8uQVnBP1lg3n+vUv1oVsEew0lpAJ8AjqNyBA7MYW8H9M4s9IxTMrK79H
twTKUYFdS6YSMmRR+JKFQwA8jTWcWnsj4WOQfcgiDFHF8U1tw3iVAWJnyp2GzDAsWBbIMP/ijja2
/QkrCsYpLOL/vmVh6K02vVYLpISIdF122teK19ICMDSbuZu9IwZ1lNxnlfLfqHfNnpncUCpjTg3B
CM4YPkhf4CCG/MBFeNuSt00eNrHzmCxodgALmyTpMPquhj0i561iIhieSk8KVAJYopyLhJ6Oc4eR
peJwix3xmjoJuh36eL1gCaQTMgFcTizHNzBpEsKXK5nRvXngJ9z1+i027TMVW0JgyWXFjHKlBQEc
bx0+ivpVzCMxSR3sxUIyIMx5/qWYvWinH1VDwf8PhXxAdhJjJesJ8eZ/qI3y0IZgTEtMvTPkpjmF
PSxxT769d+q/2cQmDQ4HTNykw9/nTMx3fZqNPeNtT2q3xnG9R3+QFCXBQT1G3PedO8qIIfZbS22y
o1v2zYI+JldgQUyjdp7oNUWsrS1+mBbCBAjN2LdicOtJ2ubv9fwwtGuHqDtYhdPAAOg4mnHvGz1q
0mwYC/JrqxfgzfgJ8CuB2FBOwVlYJ9PuXUvS7FucN6eLPKgNLoiDFW/qAvSKUVwqGYZwEvD7/xKL
1TCnNzUMDyB6PSjLY3kixaQYi7EGMwGl0HzpNOFYNk/nF7AUYnfeObBkIBNIcXpRn/TQOWEV/BhV
hLZhb4cdraDxliXkc6Sj+iyhC/AfyXZix7QRcW19nKzx2jStN5l4nn34B5RtuYjh77+39h9IvEZk
2J7YiVq9e7WEhM2kPx9Pg0kvtcewCYm49+Tng6BLfaqEk4RHGM2yj7rTVdyyFqrM2aQr8DAwrwBb
ublY7otwNMcbGYVQ5cOAahprksGmboP2mw38aW4NnBMqhcZy9igTNHd4PNoUbVLBAcj8lI+q07sa
8qeqFf7P+hWswyVGwCSjPecq+E8Rp8OiffiCBwAcfJBNhYReR0jOMKOToIGshmMVTtsrEVO4vy1B
rXRIvKR1WLr2UKNoysXL7Iuzmaenjm/M2zZOy3s49jAqNCfLDWo1MTfzibTPHETd/8IbcGOJRVUL
BFWSmavkCqwTlQDZsS5jNT1vT13e+QHFAxLnDWKCXCzD0bzkzbPIyYjp+Er0iD685qWYXVn7Qv+U
R8eq7TmBgIPVF6P7Aebv3m2nNi5+ipJCTd7rwchFrsvPhwLfTAhxcANfjdjrmkgczj0hv3hCBbIc
eRNT5wveOhMEbi5pXFIPTa8up2GiVQbrJfs38FZvWbpH44gTAb1Q3ZkQVCL01J2SFzbOX+5ys45R
2Vik7MW5ORO7CPjq/b1lSHTxOqHwqiefjDt9oD41vC/PtpiyxI9V1+6bzTcDmeVQuhpxNNHz9dsg
rQICYvtqOIr+A2InY3FPM8/acsCCWJWi8dBHZMBn/7ecRCQv8xtAZ+Q1hKPjuQ1twUa3lPGSj5Ij
W8UeskQYCnYJL3WYgLIU+RH0Dtz8kkOFDTOGjjPCRdLyuyGj5Aj405Nak2lCRuWHKSWDT+d/ln6Z
s0dKupEOkQBivp1Pslhqaq+ZVunkoe+dWah0vhm9P8t97r3gXGZyEU7UPuSPTFwjyKLVRIhVmBxn
EHJxiHNOpacgNQE0N1AuqOQ6HOIIINUVWT3mzs8ERIwKOyYL5tjKrW3dzCrEiPyYv94rQKbQ2UvA
pLGINB+FEMz9u7T1l/NUWBZwEw0tzDTgKFXZj/Dc77B4NNvC8bg0CaRKth/6XgXhB4DMFBiuqxma
zc8Ai0nR6+1YD2cT7WyOiSsvhyscub/mMju9WsKfpBRQexkph9R9GZTvlHnzMG66ALYZr62HaDRt
Lzk2aK/zz17FaVYaPb4ec/eQ09l82kjfyRAshwBSGb3ZgrTPzOjHlgxWA5Xnbg7dFp/GznG8GKr1
o4p2d+tOt6I03+nemXfpHVdP0RDDB3KFG3rx1tU4Y3uH47NmQnASXZ90HVSHVPchdConnhrkGR3g
QgHxQBvTfHmd7QtNe3pB85xj3MvMS9fazRM0t7gUY9L8rQ0F1QkR400DowtAzT343tJLLfeYH45m
dJGtib1k1XXCKoR/cuAqeQaL15ta4BgGYCFbhEKb6XIyGBiwoVFTYGF5jP3eSalDuAvQiUck994H
ri6/UPGRvr3wkY/Q1jdnJzKO1HAtANWn968ZIZOiSl5vkXIqlRKNVypMQ8QCV9olYeywjMaH2Paw
ued6nyXCHeHYki//+FLVxaWaffD2UpiPfWmqZjeZGVzr6CeZqo2Tyaogfs4AjXgom/3cFxJSf9Nc
dQiPc6yfHKJNIyrj+y7Mmn0tkxM+skwvj/ygVH0PwHOdiALJsjs3+0BZhmH/MgfzBRbSCdFdAoge
IzFPTv2a/pR9z7h9ghAxoopbMf1vedZjDL4D4I6bSiAGIIowhu2zR/MwYJvXNU8Ndv14pyCyu8j8
vTV9/KlC2c1p/aw1D51mC8XZaA5wLNG4y3LLzRggzg3NuevZGXGCLVxJUxvw/ADTw0adGq8+SJQ/
SM8M+pERPyxtD1Mv0CO9uExGzuQBPP4CNEb64jdj0Q+NMfvxl0Fdl2/wZwFaoesfGWxA1fcuK+P6
x3gJ0DMX6rB1fTHckkUo/Lgf13aMuRNUbk0KsPP92s8CWwmaTwwSYd8G9IIr8Kxt68/91t7KJRT2
YqWFgJcqqG2A18F1FM9GcvZRGbE2RcRcXMAxX+jZZ5gbCxE2gH/9ckrrbRPejt60Lo+1QovS1Int
Pisj7iXZJhAP+LovkP7/puhjz/tpeibE0OF+goT2pDvAArV9TH/g7D6RHJybjE8ahXg7JGJTjKcy
wZNy5eXMR4246/k2yQf/lybQs5Xi7Gr6VAxx4SgkuzPyvKqFUE5nBXjUFizDphEKXV/v4r/oaRt3
s4XqZN13v84oOxiIFSu031mHWNKECXNzW98YoKrCgULjZZXPq/HfpkIkRCRiyHltHRhWwQjP7v1E
0veFlR2yQYHgz4uwwxNurv2bk9i6ufnVBueOgIyngNnA3LlJTwhHjLoqdJaMNHfbS+t6BR8sGDXN
kQi3KVFMAHwMqnJzU4IGVsFNWuekLkU5qfRNkq9jsh2pvx2AWXx5oo2nAcv4OfccY1hl4UOQYLKH
euhTtBVH3tzjll0Gl5NME5YMdS26JrTOsSwNFxeWOUeJpMlzbOcY10TTHOvXSmbVxRnK4xryR3Kf
7cQ2PssoLUFbh9R5MPwGnMMLUNFnWbt3p4h2kIzRvpK7+ZMvXmTRpoQE29ox6id+0pHwQTJlqVH3
egsZkzYWEKXCX58WpOtBB1gpOt7KTdQJKKUjZ+jmseSz+uFJ2z+I5JMJngaXMJzeQ2Vxe+udhyyT
/S6ILyHg6A3ng9h5IKAYxTsrEwF3JbPJa/eh78hpDkNmI3wS4HmhD1trHl6ae64C0rX1+4Y5P+CF
av8mg0Xt8ViNoH08OUuLkln2Ff82jSTsnhoDx28iNIZ3zhq9W68V0dGO7v60GYlJBDB8QDS+DCn2
r+YWmD3Y2r3LYR18517jihjRjW+SRjAaXZL/0hWmJkHT/epkoMm4Q5ZSuxPSWKh4WlUDYYUuob8j
aNqwGxF7FeGdmKDfFKTl4DI/fSZjlQ3T8KISexj4jc+eOR+eET96jEiRLkVn7alP2F9n8puBNPXl
OUSfTSZnlJHUjI6BrtElgQrPae6RmHsXVV8sN0kKNl56tqb/ifCzXfUD/uRQR3FnCVvKIcFi3d8v
dINzv7q3dloMeJooKTmiDcghONmiEPgh5MXmWM/COPDzVy7qM+K0sGMaNYzk06kEsNyBA49+ymeW
ZX5k+7O6E0spTzPJG5/JQnJJCLuQM7wJgZEyzzYtUkMXrN6otx8NAuAAyLRPS9Q9Emz2gNIFYAXC
O2/uqxDxJfU8IgYkcKs45SxpfGzqSr2PwklZuiDmZmedu2Er8mBP4GkLtRRvlimJA8GcXzpUH/zA
GU3do0jTl3Lh79nd6FTSs2pJYABIxTeoqwfUH7Naa+bmoNsQj2IaPh0AwQN096BoGq15zXY7Brs1
vLwUXgwOSfTVPb3ozlfTHuh2sQOv4bTUKQd1z+zS6WU5AEgzjaC88FR8DTwu+uIc3I5+bLJgeI+a
AQ/G5McLhWE8T2MGx5c6mIiolGIBJOD6hyfPOehYCvF+Kk7203VKt6uwNJtDmljUzyg3evDmEkP7
xOb/tw+1Re0rOZorDMfI8glYAb+CmFXK411I5WP9XOcTulIa3fuoktp1wHUQt2vKvJUYLho3B24D
pU2FSVgRYMI5MRPyRZpJRwB0N2mP+GZJiOxzF6f2Y4de0uFN1YLPslDF9Ykpyn1rABjsF5pJ2VDX
nVFUctcLk9u8V3LZBud23AVydU+d6PJEFfq0DCmpCbZh+b5FV3iZnTU8kl6AjxC6zG2GyyDPb5pr
O1xqdLknrqa2hEjSDgYqx36Qy5L8CKtzWcOmejC0aH0TNE5Tc9ExtgkPI9sRzBiQm41NJeKDJSxo
cdjlIKeGoaoKrY9Nvluv/idc0Gc9emyIjo1dxL/rwDXn05IW9B61eezWhvnnEbrFzr0R0INEJp3o
MF0T1Uy8F5tyNJ2nFAOacRF5CSPFRNv7gcuGDm6iZatBqBgngPf3TKoQJPXABpHLcQuxBBJoPsgA
2D2sJwlvaf0IuvMR6cy0GDHiFWADyPJ6JCYZKChy5AXuzhfTp8Jl8CuYyVG7kJIff9WWX0a0Kpcv
fLgK4JMcYKeeVpvCuNmr6JVnror+aUelbFDYNb35TiXCUSE8eZ8UqlNuBI5wOoJhFMShA26PusuF
lXG1wHNgoCy2xHPUg+SWKN/h/E9ab6oRAvetBth0CEE0FNneCubqFLOUXbTm4plH42YPan9oMy+e
7nEts0PDJzhlIWGaH6JwLGNAKJjDq1vCkhqA0MdIyaCY2pUOLr76GRVpw7PJYcvy++zWdv9JLW/a
Qsigh1H6kGEenmshA+pZHeU/lVj79SjsJg0wRuw/xLzYTwFILuVX6Z9Xi1osg7xP0aTidNasvKaI
u2rBK1fgCP+Q/b/zJVbpD0ETrn9Y/K9dt8LO4BsYimGBJFPq7+z0EfPvrWg13G94AK3OKx864i7S
sC+/TL0BBLRrfL6j4VlMhEdg4zHYfBhMCqD+BSJQ6alpNKyPKtBcFhudyGILRimDVqVxOklQcYJH
ni06DDC0/DN7Hxoh4c4VxfKDyITG9ApBHMfShFHZJQDFylA87sVQYk/CraAN1EjR9+7ChLHnsDjN
8ULn2rApij1pMoyGR9J97RyVgt8OIgpyYZjB/YpAd8GVqUFH/BDnn+XPiN69fG3fvGnA4qJKSBY6
ztAtZgmM/W15TOonsHb1f9kHtACaWDp+ZNKV0rwEewwlz87k8+ygMC8/Z8EBm9z3ZT6q9aJQsd4Y
Qlx/Lmcgkj0bJtklItbVx9UunTAzv+Wq5N0g0MmuH+3WFrcoQ4s4DFpjXqVEZBpP+FXs2OnWFb/l
X02Qu0ltAbqcvLT5U5qtJLCLDYyrP6vcrknpavK3z0V/O/n8sRzH8dTgkYDI6fR2G4L+ptWLc+Cy
ghDplgKe1eOsaEUtKFMZna8ocEB6YnSJzzsor+Ao1LRHopCNOJN/Cemkxz48Zv8k4aPAUc/wS3VS
igX8KT2mvoJy/iwZQJY4cpP8D3DB0Ou4AfGg7FWZRGPgblT8HgrDVeOem952UTS8aeCCbxum5Ktc
fBDdmGukOsp67EIPasnI7KBZx2YInrNDLkNvumEQvwCtJpLzmfZsNyhGB3zdQln+geQhSNoJknvk
ESfsXM9YCRy4In6pHMhjywVo2XotP+SxMi/XDQE+uoxhjq+os3lkST6CoKafwOl+pV+lR74IrqMV
ODyoo06CaAQGC9cyfpdPYAl/zb29Wu9Zy4FCP2UcYtEwAjaCHyXwDoXi20f2PsqzooG8tcEvFV67
SC39ZMDbiA+bHZOpK2fj22mT+TTZ/SIbEcLjEsi3onTWDtJQyMnLa9W4W5lPRFsNW7A6BIsMEvt/
3uC4OqAAUELY2zSUbOLTatrLZzJ9QpXb6VZjwixSPyjHSt4rCpQ2G4lg1ibnYeZjomDcio1ySQEy
8abs8h8X3ezSUvMNmnR0y9rzlZh1Kyis0xsS3jowES0GUwCUChjp6ycZUqRs1LLHRvM7CbYiV5S9
I7S94JCrI3mH28pLj2/S4l0hqlI9n9TmBxys7IAhq98mb4UP+H1Gg6I4SJ2ncLLxAARNILdEl72U
jpA2IHgKHT0SE05tCI4bFUU+2fMbLY4ApYtJp6rZuwcbO9dFCep8cwx6FW78Oqh8i+KsrrUgitT3
+/7A+uKa3hLLBvu9AB+j1MlJOA0WwanRi0yOPQNiFv21ga0Iz7/SL+pVrn+atWysHQWwfnS64jnO
1PF2Rx4u1EFdA0NO9lbVJaDclVHILFvijUYV/oz0nUQ+3vR+U2shC9ukHzfsqOk75FwVUd2c1JZj
4yYVj3xMDw/qLrA0zhTySv+917DI3Stxbz4J1H8pwH2DB704ywynZazSYrQLK9WgZ6YbZs6vCQ3A
0ydlLbIP9aiNeu35HF+vzjfDDAy/gpA9VG2DZvHin39iOElQbc2DZ/Q/Bwk9FTeXeEjoUZosYBfG
iIwocPQkiksUOkAp9yTMPeqE8/idsV/UlvjC31jaBnBDInumxOg4V0iKf6gRXlzCeDsn64UdxWu1
71pHBhP/SIwSG9ugKDh+SY4riomnob8RFLgNJaMBfRO5KjQAriy2tw4I+ajLuHAMGcyZq6LqAkuD
9Mtyt4PB3PnoaET2UKuNoXnNOG2xzMuwb4ybCeqYcH9C/JNKLnd2ZFcZET1+H11WnF8n5egpEB6e
J3FL6YF7Ir7Jv4+eWpO4QqCA7E+xbgSfv1ynoWjOuXKWwliKN6eGgpU5s5OyTLZDMcHKWhuO2fZI
D+C+J9u1GhK9vnBve7T7/zXo/MyhkgmZpCyBmOkM4xvvfplhCpbi+FOD4k5Cnss9rEnAAvuBS1au
APOl0LPXMjdomwuatPo+/qd16vX9bDd73V1uzioQ2W1UuWOnaK9LihItEmmWHaOlW3Rjj79gqaxc
ImToqJHcjhvlnOMYUUBWXsl4HnhgIgqeCwjn1JYZo0HHJXERyuyEpeel/yzFT6lSrJptEIfcNvUq
BoKtC1ZnEpxR8mgRe1jiVOFDOX5rOqY4nN/70zJLmJnQMWdHAnEnxdf4DE1gAmWJoz9vyZb1aZT8
ugA/rgGs4xhi6eGY/09iLoMd5npKSnkoMWd1zebeFniP7e+ewx/YzW67cG7FGV23u2wXuaxxEHY2
HOZYKReHs8evt1stErLeQJ1E6QutCv+7PEaAm6Vscxd4q8U5fLwPG5hZ60Kb8A4Wc5n9///fGexT
w1HeElZnOd/gZKeti8H1qRSY1DtW5VSbqAo3an93rhYCGaN/+bCkqS8ZhebKkf4wEliUOEOhZEFX
DxkTrrWK9Z5QDTPe0yu3a5YOnxbVpr+LmbLs+6lMhA9mH0we95DFveeMvHhJnm1P+SwbcX2dnaBg
rl5Dyx5QyZjulpfC0c36lu4zhqE2VUayY1H3SMQMFe0oZy3VVRHcbpbEeGeQjgxGbZy43/5mtDLH
VT9VXXQ72RyCxJdxGpQfwlKbwCSjIm1lUJLA4PSuibdbH6t85w75rlYsNlHTUBduiKZHWuPdB0os
gU+Vm3uAv+5drLUIo27a4NbJg5VhreNsbDCQ1vaTzusR6ZST6uBpa+uZ7J/80X003P2ymjhLqLCK
BaZfvokYucj0SJaGxr4bB+rwtk8SK14Yt0rSivUPUjlc7pgZd8oJg32tIXKayf3HC8LK+z1fvK9R
ZOLj8Kt6KVXn8dGipq4s6djmYkMJjDMSGYNPuqvqRLCaQvWHQSCkf3TDC0HpEiF+6CjFx8EjV5+u
dV6bV7p6R4vYH7W2XCpV5gzndDgxlUUt/Ucy57nq+QiueRjE9c7ziHlNnGe4xYdsrgeTWlciHdBm
uFV50PwDINklKCwb1zGPkCwUPeVlrIEgfbCli+uRfda4ZZcyy+5SeugXwa9a1wbmTmiXzq6x3erU
YDjeaxZcGlwOxGcLBC/DkMEFA6iQdy8j0ApfxNKyfXNrtOL/N9cl5ELXNx/UnNgUHTfv6LI9GtCY
aDiMRu6oazHvijTLdCd1+9qcs8Y9ZXLBj0QhTsWoF5wIwSgAtgYxFbQXaWC9EO/Y2Vk5r2FEob9h
glG0z+RGGCobaDTxAtviYknztQnqGGSoqdhf+2czdR+sW84sbT38dsMNSZMXvDnY66Qf+SfjY2CY
3lu50hsFXtT34tX/uHkDJQSGiAW9ZFQMO3Eba4hrV1RSVeflkFg9rmVlH/0bw16eJgyrPTNnswsH
daNZoBBbG/ZwetHrYHwqu2gIiW/sy28qflGCTl0hlULRIYQulafR/GTSrMN8ITFHBUO11M+L1CfZ
qCRzPzGv+dy234MrY87PvpkJ5gxQWoduSZumbTVA282pGC/fzMMUTYVzs/3r/i/7H8mULP4uQ5Ij
94nenW9nKKmg0A3taoVRafvOd+6rDG/tiRNN3E/zq+dOVVQTsS+jXGA6pWHjIQx1sqCldzX+IWXP
Pti0Kh5+qTN7bu+s98f/LtZvhRbAHUJ9HVUR5ZuWdXTsApS/+I4+OJlyDikhU4iOTWqzR7cUrsci
KPybEtU21ICrFyGIB73c4hqByNI9w6TD3PAfKHvOSAlVk9voKkAV3LnPC0N62kpp01kXNib0aA5/
t1/iIM97qvkwHu4lZi7zghAOLeAEfXub8r7mkektSiOQ4MSQR1WWYhBY+0bH1QRrzU6rayax8Pg+
RrwGKeZ0ZtDstWvdgrpF4VHq8RtTN4AJq+LZmMmoRqVKBZxCMRj8K0TYeZuZKSZdpTSuJLlr/mRt
g5fbsqAp3TSYT9ZAHRXH9dZv+QlNV9WkJqTfzsKtQkqdqFpPwEJnZCwJM7zDbwJaWnmKqyT2YIwg
5neVt9UX3/jyNlryrCse8lkl4TJ1MggYplhttxM1JsVsuaZLikWfmlYcx2UenNKx6MAYDRuqbXcK
GDKmhW5bIVm2J+J7p4FyDtdAAmsCp7HWJq6+SduxjWqJtJJ9A/IeeTnX2cuN8YFQ1+mm/G02hOl8
d1H3ddw+I3Cm+Af5Ea7a+w9vdTC9m0fx/Bx0+1fZmlq/AnBYnDIudacBz+ygH2GPd+oxge0/LceH
1evq3lzavL6j/geTttgiwR3KAT5x6RkEZIYMRtNzLa7u4iZugXQhgynAJlqrfpdGOFlvAG/8iNTU
v79OxYko1v+gK+nBy6Se5CZ5E5vDWqgkP2AY4Af+ZWYowLq/FgEtvEWMBPkJ9RBtK7kwnjWAQmL9
z/SHQZYlla/suh148eoM9uGVTw6haRdmTsetLIJ0S2K7Xi82pDPb/wQwbDKpF7RWevpJj7cpoQup
Cr/27Ostf2weXx0UPzvngrHHeMLBPqcMLdsHPSDyaj0TB4y0NUS5cVssgWvd2Q4vSvU7bQnnmN14
pYolClYKNSe1g25N8c3uDP6UVUQPnD6bY8S+gJoU6Ri+/97vKjbxO6ygVb3YGitbuYOqGjrAVlEz
SZmJPXvcUeSDNiXGBkjaibEq9BPY+fTVz0AOzItb0wZS+7YVlcFY0ktcXj1i+AiF2MaNcbx34v5R
qgoDvvoItZnlO1Tuixd694XcrAiu+jGOaf4O3brNeYZqu2XiK7eHCcTvQ4CBeU763aKpPZKcKrlf
XUZp620TxnzED8OVZ25sSy2ysO6JkNczINQE6d7w8f3S0cj0UP8HX7jtq+uFgp4HYVo8i++ggcR1
g3g5upxIQvQmujYXRnj0vdDgV54DwarbHZDW48+ZJEeNW9pTwWKngjELFYw/THXg8tu/bTlXLukD
D51bCp8PW49YFaa97DGfvt52isOk7wBIjkmz1qEqMagnQazpi6g0VrWIxYY8rSQ/PxDGUAWySu2v
FsxHloHRKAclxmku28Ode51//7L7SftNludRUPzuT68AI+p0PMwGdC71eeBn1Wqh3+Sal27wpqzd
FmUHvg5O9anO+GIu+RQsvcBqg/sWqG+3or2KIZqofdnUgQVY6uugh+TFMLM0OpYp3YXeMvCSBeH7
UmEpfjaxP6aK+i0ZDPIiiLlEpc8tTALdxPu5VWQDn+zMYxbV/W0nAToZ+Xt92HcTGXBypZug/63T
PQQPq4c8qhDnLpmjQQJx0k7i095ZZKHuKEwE7DN0Z0FPkGL28YBBDSaaHUvDBuR7hjru568ha15h
CpIglw4QKtEJEVuHDonz0Pna5MPOT1tSUv0OFc66m9jw+8/wYUTvyiNQ5R9NZ33hOiH+N9IBh0+F
A+MSJ9EljGahO03N8Gngs3cEfTU0d9/xQnfFZPUsKkjeMVv5snkLQZA3QVXywmq9jAQr8mYs3e4s
OVPHSHrkOU9nfmoY+wM0fa+QSZgDS7xvXcGmE/YCGRRb313cYrzKJq94UDBHMk0LhVx4eY33VOmo
fvwyUuF9YbS/+LncA07GSApsZHyo76lvyIb99S3RUna5vB3sZFuKa3nRFoqJ/BXfuXuPJ4+CznrQ
ZejNo6vWUfiJiiJQXyHIDISGyjAKBMcMAeXAe3DczaDPwMeXodo4QFxfKRO07FcopgcvpedxUY8d
HZyemtIL03njK3hElYZdRnN73ThFV8p2pn+9MDeMo3JiMmbsg4An5QFpUMDqNUAJIFzkuXQ3IRlH
JD4v0rxPueLQwAAu7MZKzgDa67ySP3zs9w/4KJdIKc8Eg8HrkCjFi2jKvROy3fQUHqgrd+7fS/9J
LfZkceiGfVd/G94UHJP/KHj9O2Re5pC5DQkmd4TSnNpCmsnSgzLVgDrgml5PVpluRcHR98kDua/a
aH/95ASr3yAmGB30ZsXG0M0PyOUfXfCp7ZWcKPk8b/g/wSZfn+tYPRNoEPQ8W/lBUDzCPRhmr5BJ
0Rtz6Bs00jKWv9li4qwAkGdM0G0d9MIKtexE3TCu/veg28wMrVVup7QQNKC1Mp0DITjlz/CHtRPq
s94qhyl/mDoTjgYdqEhnC6CSQbY1d1s0/6Egzl9q1Btlvwa+WbtNiIdFi4XqA0bEYv4wQfYWFxWO
gmxHo+fEhsyb8Ndo25YkUk3UINfbjA5a54IZUatm1SnAc3MXYm+gAP7iQ6qtAxDcGKllmMGfLqfX
iuvGqXz11rJyk75ikSNMnCMedQas6USqVTisEwTOKR58b31K4ft0MYaDQwVvRIetJMLwuUA+ZAF6
xZ3Fbec6e8UJkCHYKvBoP11cJY/dg1hw749BvWK8k9EUCW1NGeTRdFhW8Z/W+s6SAOWC+kqDyW6H
rhdCfunurhupcc0VeT65fHMpKNEc6SR6BzfRWARCw8dTVh9tz8oBLvUNrly4AV0Vdj9rXESnixHD
gVITofCOAZBoa/u853ePydCF4pZmYDYLavvzFE5oNhU4WynTKhg7YqoUIx5Yp7sg24AbzNqNsHum
Z+Eny2U75Q+SBeAQfsn5XrKIq4PFclCWTNvw45z7I/bcXGT6QT5/RiKuNcaUQ1xEH5SfgS8ibpTp
mFx+cWUm8UqBbOhnrye+vf1nfVmG1sjMNkuMZBAyD3gPdIvawBtLFnVlCDIxQ5LJs5yOAy2KHiB2
QacSY/RFgCxsg9KSRlmj0Na4iNtFwMT54sc5tTxIV1VG6rFBVyLFItNs3wXsfp/ZuyETe3lv5qt8
kmaQci8WLuKdasmh7ywyAIsN7Ab6K9z7F5ahoJQ1M6+XVEJo/7BPOhsYvSg+IGslaFwLVbDndZjL
lsGi30RiGx+hY373qzjDq63DMcX3eLPXoe4mx6vDvehubSr51tOnrITMuuJ/spMF6BAIeQLoaimF
7SNizOj40fvAFe5tCSKvh4x+BCbzRZfFJ9csTA9ncQCdNF/BGeR9FkxiwybgbFc/iOIHsOUrPY2S
DdOoLeQcl7h7T3rgY5dNGBLQaRdmgEbfcGB+QoFj2J2XGqjaayolPt8c+KhfIeGrwS4Dmb6SXilh
slDD+ztNxrZ34mVJhzTIwy09ZoMTzKiKRuvROIW4A9IbkGt/Wgy2bSclxYKoPKZlxU8AjQhoQ1OU
lshugnlQneJB7b6ZfOMteZL9iNsgL7snsihuLs2RDJP0qZgImIYIdbkE5scyQ/FGAB+ZoKMzwC8C
zG+VeMWexCfa9BMqifi0H7kLAiGRTRP/SuYfIWC5IPGPn+9yxEz2HqWhMmBt450ApoTBRdMjtFta
6VJpSkiaiOaSf96ipvsbR2HzZ42RwXmBDuBbmmW82WZRoMeLFGXAI/FxmSvq209PuR+jtA9epyaK
1mfQjlOejq5QmunX3vXKYC8eQqKIRlqW8Hvi6If5Fh2kCUUHEzq9FgJJzPA/+PALTgQI0oIVLu7Q
L0Slxg8j0IMH3f4o8GXsc8eP68FxqngWnO1xForFfFeesHf6NSBRwEsscN2rjIsyXk0dyUk6S/G3
wh4h6fuiOlc+rQ1tcJSe8LE3fWcxsahwuEiFT+npFoRA29PEZN6v7nZEgogLkHxFNi388YanukUB
Jh2krGFb5sPEO9+e4ne7TCeHxD5HmNv5oVfPl4Y1gu+sbLbUU83B0U8ndB0TZNSW3rl4VvyhF4hL
nuQWqtKvOFy6UbjU9icOH6/Y7vc/NggOPIFes4c5uzEDZnA/8cX6FmvAoTrF/2jS8Yeaxp9x4Xx/
o5l1wB+O6CCdRDeFeah2hipWFw0DDDTzqH/2zaZxQegItm1PW8ryTlUslQ9bYJaYEbPV+kPWThdy
u2JrUHdS0sfaeIafbqCA0jV45qZDIKP7DuOaEqPQoO5Kx38OhK4vDs/1hAW7fpaTxr2nI/Nw+fbJ
i5+71UfMqEECX7TEjNaw6i2H3df5QNfmmqz/AlV6AWmjqrmJ35IuaFMyfWR786wZcFg5AQdW8uLF
UqjGYciPEI/c/NFy/Boimsytx6ewe7L+sQG23Rw94bpFceMmJ7IBhb7bcUuC1cGRaWugHFWLq9NX
itkyGdqC2dz0fx5JhtxahP1FL+xK+XtcPgbuCMLI/uBIZMpl8b/0jYHUno57T60a/mZ1nBIqh9+W
7jfBQ6fQrS8fKn0rMf7y4/yV8yRHl2wBq6ZeT4z/3jBpZK85raMp7U9PF9nFrLac+WO8lPIPAz0k
GYZtk/i9TTDYeDdhiuUE0PFthr9pGuKY0jU0tGeHcSHNCSxoF5cwT1guu9Jr9SCK+RCiBg4xHsxp
+Lf9jwLUNPFAZmg4UbBsmDCLV3WThVWTb7LVIdcJlvu4Losh3y7F5mUYg0TRPReDthOMuP9rN7U6
Q5VL/muI7udV6oyXlOACowgA60euY2jlIuQJBk5IBDHLmxWi/I8QoxsmNXM1bGfyAdlRtl8N9Fvx
ARz5XBI/Tp99d5A5FEiQB0AThcKo5s8Fr9qBZA0bQX+C0at+6acy8C5Cv1ppRG/CTHWQR1nILLGe
Krr4B9TSPjRJxu+BhuRPOIRVD1grJ1jqTAUtHEnfW3TyPnacnAOwR0vyNSa4NT+eZw3rQTKNVh3o
vV5xgfWHR5/SuDxvBKPWB0RqlU2luPhPtS7yTMHWvJPZNzOYYylE/NInR8a3XV6hoPHzcbtbuLcR
6XwBQZ8bxAM3rLRJ8OT0jicreShBqdeiY2zrYvX2fWjqe3Zgn3og1SggnDSdsow6d8n5yew7SiL1
P7K8Do9WRYjh9DOR723N+bV6M/4GqbPFmHB0GeaCi9zOMJf98B3pk6dD6IOH8werWasxJwnAiwXR
/hFKvj0C8Gsm5I+kCy2v2zZtxPHAmgztDGK0vYo9wy5sacczatVgidHvtkj+PewaDooocpNN6Dqf
7PgOkM0ZKqzGsEswiK9dSaE7jBz1Vlbj0bZUooTSGXkvk45ruresL0lp3B2/a8CHImddN2YGqcXa
tHD37yiq8z7ZJD8ZxmI++BVfArlm5fBfdK1yQuZKMiuaMVGFVTUF8dPey6YQon05tCH0bBFhtfUs
7XtsMwOwCn+hwESeV0Eip+6fennPLtv6fok7gfsKGkrHPZrDYJZnHUF8e7mn26x4gae0FHVD3VHL
U4NViQAUCPtyx6J5nqXgOSGX1Qfpgch5wIcVuXZFH+MXUUZFzQpeOSH6/d0Ckyn4A1f+MWxYwHGf
nEH0otoc/ItZakZXH//cBdhe2JuhRt6RY6RyFhfjiDLmuDfJfzRp/SaeYF5tAwBokHTJel0dK2Vk
NH7P5Lm1JUC4hbBY+0231N4GyKkn6U3esj8vvTZU5yzonJ0Lh+kyKtxcFvCqUBpCJaFqBAOuz0YP
EpN076qaqJnza2dWa/x1PZnvVco7nlG82ShOeOJERuDtd0+xuTp4TT2rAciIu2BzmFQunzrC/eTt
YIYP3Unj0JMLL83E0MKqTMh7pC8JNr1TOMamAwkxM0vJms6Gwc+UFucYIUAD6NMGxDTA5KUImvIX
0IDMxU7kGLMqNvtycudrWgzFqfyLhp38lNjzsBUNXdllQOueO+/1Wop6BuFrWv7as7znesHBnDHO
DMXY2bC3Pi6e2b0SLFTn8zkvI/rcSnxLpwlBX1AqGox84tO2kSneSZZD8caJ7XHWYZmrlRdCENwE
YrP09Yz8bw0MuMkLHmegkW9yzeNT+JIdv25OBp0xcilvtRPClpAtLqAtQl0GG9Er9li3PXv+xcE2
WtFi5oVtecIHQswU+FaUicnV3UJe1+g7f8UxePucAGmaIcNw9q6XaRX6+kgogODQ+TPhgKSI23Ew
zpXnZdJtE8VhGEUSV88L9fb7gOk3Wk89fhkEuIT361AUUNBx8CNVUwbQmjcV8cwt1D8m3rs1+edk
P+/aI/owvUKUfdsdRSQoC7+kDwsPpafG0l8sgLM/YabukHvOvJ3R9A4btpice5ToEXmtp7G14Yn5
Spd6xXD9ZgCEjPxBQ8mlPtn5VQHDmwpwFDSCHPYxzlxMrkH5VsLXjPHG+1gHM6nfF7bBYOW0Q96f
Tq8AOyKTu0uX0pF+JH1jzdgrLtllWOMXbOLPbiCXQGYYvGBqp+lEx9yi2pBTCUfNZcloC/sPVk7w
KYw+mTC26W/jJs7T6SHKK4zaZey26nEw/4scuYZ+gmBMALkJa0ly14+/IAWSuFzBdatzF2cWSKvO
PnMaif7p6/fei+041kHyz9e9kQKCiY63hmEumDir0rKwoY/ifteyOXa41esVDZlOVF5YZM2GfTkM
CCrwto9J7IsWIV2IcyVclVFVbdkNldBMnbq4klDgEel5Bm4b97sgI/BG+OdHM6sPaURiAtIewQIx
NozQdAknFMBtsuuAMg0q0Ho5qbWebV+6OXZ4UeMvH7Ca5qaylL8wNxfvje0DmJzvdwJ6I0OROH8z
vvYP0AQXZ44Q4ELy68DPHs7kQka/2dtiHCa7KGIovRtqBboTLxdVxVCJh0URGmZGYcvXl/1CVIB5
PNtNLmyQ2Rm+yrlosEJNNqmRzErzrKxaSdWU2bCSkj+6wyNZr8XynirHhPcOOxmqAFK4LmD9HJdq
nMD0tCh0FrDCGkmfAwZTsWWzIoWgrD+0iLb/EIOltZPHyqCS7mC4ogIRW6i//K1EbUls4LZcoIjd
YwtQEo42fjycCSAsCy2l36cOPdEpCPtF3cDbXtyr6A2zSM9ALJ2D3zSuEAxgMOhheaWcBuQUl/HI
PIFYwNJphGane6c4wNBQ37PPVs1jayQ7tQz+K7pDEW855lMal6POW+FNiVVZYvQ3pte+QSqGVuxB
tVEkefA91/M9Q45CQqedgvvLGyh0qQrDe4igJKSlZZYTrCA2KBJpIeLwKSSXQWL7IFXHZQbXSz4G
8Zx8BBviUvLnAPqAGisaDbv2FmTuUEIG7gplOOMaQJZkUQ4vyRdCZ8RN7iHNxUTzcL+d6JTIzCHM
QUfROLnhScyhM9G6IVHPWFCPMpg9A8Oz724LjaASi3o8CjCmaPUpggxzA2S8TLUl83V92inKI1Wx
fyBON3ZdFRzqhVRMmyJYFd1Vgw0fJfT7eaHdGF+UgFiqIlVbO2v9sstGqPan5yphCS1NPv4qAgnr
Wknw3OAGkgNeeLFhz/ohbUTyXret8Rpy99onPkFbeLG/N3qS8AhQD7QIzRWpDU2dbz5NBJ3E19DA
as+ek/LiSExqNH1YuYcRtHZQ84t7Ke/iX6N2mPZESsNMJ5SwRWEfskRTcI3K4VMutE3/pp2rk6J+
3+7UcrPi4wfXPQ1uXa1S06qx+CVY8zeuqIevUXwPpnDHrzBd2o2GBuF/w3vzl1WCggfKLaHtNvXU
dDb5p3x8gk8Pz+UxeGI4MfoTuFFAGXSWeMBSycMu5uEVYPugWgOC2CK0Y51f/F4f1zw35G60z03V
McG2t8O/XTGuwRNlvKB+c4pJPYqNfgLc+k6f41mqF+TOLEKfUhSxiDm/DisxklPMfU3j7mlTqNd5
D3mjMS6Ywtj+mjOWzu6R5nYQdfmfrABUtr5A6R5AdhBKNYzXF/aTeLXg5eR9crS/9iUUk5QO5P/z
NXMXyOi3BIBA51ihDbBTFK4feZjwGgPDAPX+xzgtL62iEOnFFOnY39k1hCAw8XpbycOuJohGzXfu
n97eiHUorfdC8jkbwmVPARhZ0+30VZiWNjhntWdaQJFKQlPQJb/QnzqEb1EaAAegX8QqgmWAj61N
K6mYZaW2HO0ibYHGCcPrWYSX7BHwWzj9H1kel3Gojv+9D39hZtdymHbcGw854h0uItwbIaAyatXY
IBtOMAl1XdzXs13yqX1S56WWdNbI9ChGHOVqhbXdZ+XER14+TwkcRCCwycO7d+/KdkipsbE3tgc0
mjdzHiAuKQyPlR6nZV4gBVt1U0UWhx5eaVImGH6TFjXZldRotuorYzeeXcuA7CPZJyRRHDmRy5cf
1w0DliKOxbMWM6J834vII7DBUZNrDNyF1TKbsPgGkrt+W0EvrzFqrRv0GxaWyXDe0pltM34x0NRy
Fw9BjXXyukZhkopKqFgT3WijMHZ+gdxv69AYin2wQlEikT/sGI+i6T9JUWLyjxuytTQOsAGj5hBJ
i5uEki+5+06w5qsD92gs+u3Vp6bNWn6Jiy6E0JIQzcQh1r176sG7bWmezOTiHiFc60x/f19oYaED
i/fy1WrTAYNmYELqvinJ8HNwliyW3Sj6JnrUF3yeiBbHy5G7Y1c7NYC7zJFPJ+eq6/3VHRu31K4M
56kGYVzVNYxSJM/5txNJ//rN+501NfTmiZrkvr4R3CclggU0IMhAjjQlcSFgf0mYp/DgtebZnB0u
TaOa1traqep8gAGNZPmWuk3ol0ioA3as5uyhTZaZu1Ic8mOogLd78jSpf4J8SlEj2kEm/kkYLMz7
D44PscK9OJEx48F0cx9WrvtS0K0sTS3Oxl9xwKw50Pm2+O/fTaSW0FCN2bnwvT0GwI1lAsxoBffg
gG7e3x6WOGmFTtK0aOebd/H7R6bQtoD3/RwCCCw8WFoefOhJclMCAkDaFfJ+repbdShy3toOgXd9
uspJNlh12cbZgBxBtGUSbOdMTIR2RKbCcmBowIhy0JRVQCB4b+SLEtmmokFqqI1g8C8TiQYqJOWf
LU0n8pDszsCfKewJ1dOh0UIUEMTTbXeRNB3sR9hGDWd9ulmYGCPyAwfeM5HCPM48XUuxW/xT305+
flGyzFJBvmJJZKvTYSBcfmasrC5bDpijGPxaPvLuzJnjj7bhCQAt+FQZ0wdmjmUkXY414OOzvfmp
2o+R4A3gcQQxoN3SFmxQSUYnP28T4yiOcKAYTkq7yE2isf26bfcgEJ4o3UnI9WOnPkb/ESpW3fpP
mIWsTOHYGbNzB9JLF3FD1/AONgJmLU89xidJn8WEEVKnfpa7s0xK1YkoS9gdeKy10etUHv7i5CYt
BIp9PDl+WtxtTGPqPQlOJQUVUmBL7+Cs7+lRG7SsQy/aTujX0oT1O8v/6A3vdLoI1dnSoVhZyu9j
UWXsoF7fSv1hHnJ3xwyTvBBOLGFgcDLgxICi1r1JoCut3uKtxuPhicKCd2RkswRJkl/zssvQw2Eb
qKiV/8XdY5FXKbXQ59kspV5HClOIvSm9EVygzK5zgCwkZibRKKpHaGAU+XRnm0DvUOyvcp2esKve
rU1/7gJajxQig036f92l47snXgdo/Y6WhOUtrw9BVmaM+Kdvvz5S44iA6gaTgMOEb2+rb6kWx+jS
XumoY7toM6c6Ldt513JVZHVftO4NVznls0jCMpckMHEEnVGk6R2b9f4zaUbq8ooKdX+CHRphX+hm
+UCURDRjGInPQ9l3bmzPP+thF1pRNtPp//9cTv4mJ2/9ZyMUdws0CiuNKogXdHKp16YHuXtgZ6mo
fqm3QndzAoqB7yM7rOlf8aQLFFi4wFFi7SKWu03tyftPL7VQ7Cpfk17VCQWkQu5jxLzP5q2itUlB
EgC9W2IaZKAoW1m6va3YLZ4CT+ckFb74ZjIbBGHs6G5flQvGdxlx0FYrPCj+9peLoEltrvfMvGQc
x+wEwxrewdPiQsq1OwTgquEEBOBuhiE4reNcribgfdFpcRSXkeXW6jbR96vz8gxUAOHMKgf756qf
3DtP7snYVm1WQGtBGWYLauSR+Q4Fbidknv7Qba9Ac1Hw65x2mLw9i+lAwav3OsCYUSTL1Hn+wNtw
APvlG5f6Qr7GaagCS0qybFBsQ/bvB0VyNh3PeuY0kkSqEAVQRyCPoSao6jrJPg2+szdoA3Kk6MQi
7Ar138yrbUD+Lsb5z4WMDCp+3ZCVTymz8YbPGJLtiLZ2PxcNH7Icj3g60XF7zEm/rQvYzEDcS7W1
2NsHDSuF7+jQqS80bJgp3lcx1UvGqAxHFBoNmRoMWaBWfnO2cqkL2vK3975DNBQlmfcY4jDm2pcn
/onLNM5BtpdFyQOHfgcWaEF+L8cZZbSfKLA/uBmFvE1hkiOu+uiYuQ7918wqKYDicAVkGHcDqalz
7ychtNt/2EwhT/BSzfYkAIsJLM2dBxI6ngl+xU3NFZ5zdSVV45x6p9WqkOGuRphZMVnOfDgnCYNh
t0ngbvk833QfKb2AB0uOIrECwq4zwP/f9PL3AlUX7YKcqqOKKyONs9RJOy/7CuPtULPfCefHRgBW
z4WC9C1p7GczXqvPTqMY5uEkbfm98oK09Qu7JqryESSYAQeWsLxsNV7kcEbdMeYkM2Q7CMk22LqI
GWrqr3ZPmLhBa0/0c8kGhKl4oCiZwOEQLYmdyvX10SEqjl+3mOlYsl380yBaGmziGejWtxYZfTun
2kOPa+64noNWv0Lwe0aGuvGoLKCaXUG4PlAKekDyfYDHO0X9Vs22zbSbSY+6/krxJ2gUXZ8LoFKM
1akFQd3ic1d11QszMjbuVfEj+qoFrwJGzYVvfFhJu2QRKwuUVy/lvlXr9q2ViFWA7GCQ1xfDbmCY
jl4RWN3AQ7NTR5q1tvyhpzXrv3w2KiYx1IADvI9T2qPtAZvCO2kUJwrpu65D58oLJ2WKu/pasalA
5LxCKF+08xZfIIaCFla67sO79IFp1ovk/33Y2lTaojOKM3NlDfsIs1KCBr+zvn06TY78UMwdqyak
CbMlABqQbkpfJd63SpsQ3OQAbHWczULKoVMLx61ntbsMb2qN+uf5KnC9Zb20b8jtfJpqPhxi1Beg
MlbrTHJ5qWtBuJoelPfdFZy10eA1gl3ddcuNR1sLtNWBenfR+qClI+Uxfzo7Ocad6r/12M9MWKvZ
Xwfg8O2KVmstqWzpebLpk5ahq/QRt2ieiWNAeF0Eq5k93Qe0YHqMjHwql+ZrTxs7sEKYCjqV67iB
/oDUIvG9AS4BGcXgd+x+K8OCenLntWkB3RydqzJt9xjuVRrAPMeFhFCpc1RZ6rnoi6f4+IWKcY8Y
V1qiaYiLmZXG6KQRz0de4IFHEW9RmO4y3+yveX3ll5BID5JyzKaT4JdpoPX1doWu0lwNnYrfZlq7
k7ncpicabPqIMGxQ6m6rsjZ01cqntXA+jFOOgcXVk/+bYGOM0XzVTQaf5v3IGCEh+M+m3emvI6UJ
OyfGDvjj/LVHuCCr5sny6uCfKv0vr0mk6eCDeHkF7DIAcctpX8RcMzswOg2fFFES/HjCVm32XCC4
xwtOFMZiiwPMHJDnIyjDkMG5WL3sU51RkH6WkbyyYZSMrk/KUrYcGXWfEOhCP6AusPqJePecftR9
UhR9Y6WXv3TtMFutDmJppr7meTNUKNSMzsEMHgwv38tsMsZJiDKiUsnmemnsP84jgvw1zlBb9ccX
TenAe/sfTo+h3ZMbbtbEyjQXZ/SApxdrCdmbAofdb5v6l1cFdyuEvj2p49yl2GZp+aAKtaLdNXqZ
rV4BWZig6KGOhkCTjfKsRsHXMtXClp/Shia2WR3YgYJg66HtOZ6OPuRdY9PQKvfzjxyYNytA3KIm
otvI0SM5+rzQwv06qBGEqK1BNIRqfTxDorx+dMTV7kO7Z71WzXEKFxDC0Jn4KMVrDjHjcwBAp9yp
/+StFyjwJ0HSnExdGrE4bK1fs38dHeVY7MUto3vBBrUZhg+hr9vFHPQz/bZ44irR+E3KbysQussn
Shlv4BVv+gIwdHwxY46zwjiUJyMI/HKnKPeJQYU+pID2QLr6e8YFP82ETECLdX5uiAXvGymog8sF
Wv0cYBa7QEUAwBUOrwSvRIp19KA+r/Y3QJQ2en71IF7krnmu42QeoHu8K19xIWB3bZDQz863Reni
1HuDsesu1Zfat781TbaUfrZ8jsY2eGNTYOpSDcXPBNWge67fxzP60rOkCL0rumcX7rolhh/2f/dt
DuAy+0eLmipZQYDodZYlaT0KF2cQ4PygFNoQ5pVd7b/rLUJSNi2NkmhzYMAB84meFvDKt1eUexmJ
dpOE/GctaDmssOfOrtN+sU5tuqHSjG/a7nvrC4qe2G9566jK3tKtJmGTYr/YXBkgLXAKyMXqCrnt
ZFZyAf1QbDQTI2XGrWcj5cJttkq9hOdwP9zgchnepRicSKNgo7a1zGwY4rj7beCpXPIQaRjOg9uG
ORwAmnMVYZHxhsD/liVszET8aKx6jw5mB7UV5EFAsrO3mrhc/KB5ujk3dCqv+17HIFJ5NfeXBTKm
MNZwPt9Q/sf3l54XNVdNZS/IqT7qX59BT0VRPN8NQzc/sTaw6EHz5NW+NpfefoahzU4HV/qXNGgS
vtiv+TJ3s9Y504lLpJP9+i1itHiDLWlAroV3mFz4YT9IQkIgl8Mm/3vJnzVW8BEwp060pph6rGf4
uaibwbXnM1p+wzwNYa+K4QZnRanBMaAa20DBVTOfUflWwlCt61t03GI3BogjasuZWUgqk7GAAqNA
Pm+IdtBBfdKL6O6YFk280juP8BicVXpfeLH8DVWLsQ/NUZ6mFh/GfTcSoPFluR+YNyF+6XAS6vtl
ckkhtijb0wrS9W08wuKq6j9eJmsYw2XBNhAg2miZftwsX/FP57wOCEjtD0kRtk5UpsOMag7/aVTe
kQnBAFcmvnmw188+TnQOJQtRQfQzLbM9YvNuTjTOSbT/ODoJgCbtsmebEKvdPQ2eVlBa+zH5IdqA
byecE5Bc26Alcb6qtdwHwaP5u1GnyjbhbU9mtN6xOYOpzX2WOB35RcloJpz+2Lo0JVLSx8p3Du6/
J4vZvF2cVikWESDkvKYI1i+XWJIxEzA9RrCv7IGxpEYkw+VCSbWCx/51tMCVEiIknbY/gGUPShgZ
HUoK0VYGX2ruiE2wtHBPb8Hwtywnj3VKx1Q49Q32tUaxoA+4v3MijZekbcxKVImxPWIy/3wkfNOI
3OuwtPv0yKG6LguF3JUbOOqTwg6a4YMr/XCO02ELzUL+3kq+fTFMDj9OiXKN6/6DF5MGWvTKoGHU
KaYu8RyxSReUT0mUpau4/v23cE3jDpZC2BgZEc92Dzf1gZBCcM1Q0weCo2nTPoNYXudbOVNfLxw+
rOoeXPj9DxuFs4n/B22ebAOMRbKHqpxkeybST2em7NMfM41+3ogD2I60fKb54quTLdOQ4tpwh5is
3xqGC+q4kMHEU6U2IOHZla91r75by9v9P/4PlwbgG7EBcD6UTV/ZRBjOAqyNiTLfiItMnsUmoU6O
7zYrc4HmP81dvtekuRKopFb9ThcxWNdkw3u/o95JaS2VKDTL92erys9WRQnVZJ7FuDTQY9e+RW5N
gsF/gBiiuE3qoDJvnbU8U55WlyyhTV9twCclJ7DA+BUf9lRqt/nT/YudhtYL5j5iY/YeQplgGApH
OkhABBc5/5fpFnJUSgJUU7k7cfPAQi3i2YtxDBd19ZC3YS80Dma4eCMEQxaEHgs5SpDbqZIe82US
o33BDA2w2ERnCaNa0Kmk8hsZcpCWXkovA1Y5pNl+klCymlJJP1oebUzW4PlB2az7yCm7rLK2zoNc
TNCf6AiILF4UHVEsUCh7wignNveWXONql+2aQ7eZh6d68/eMkBdm1lIZVLic86c51z6/Hkrk7Jjv
LEpBIz2R8LIn3lDHT/fNEHJPMaQpOwKaE7Dn9UNq2lpcVUe9pEBVocuwdDLtL6i4qpnRFi7z5BUl
Ykl/z5omXMKBiqHZJzsXwPiIIEPnZRx5UeCEsDuNWV5ZAUbMxEAw0amomn0zJGgvwIAsQmqmPHGd
UI0CIAx5DUXAJYU0b4yDHFFGVa8UOwmJtGJW+Dn4Pey4/ybwhsd/tF1IOewSNvOC7ktEiXFbWWEu
Rmu/LeVde0Oxdy9z3OUZ/AYZn9XhpV0MWDjlIs2xlKrIIVZEdJkbn/uGv86V+kwSIrnooHwgkpFB
8WnPXGEGdEC64BWpFKyB9pVT68UxwDEfuowFoZIX5MdJTEyBL70KF+CRrM9oLlssYMfLmx2XjlVm
uNXs1A2vIpSIdrGjuluXJ0NS9EtdvCCf3esfVgxNrSS4cJLDtEPVrabgjTv9xPO/RYT65T5WVG2t
NpOsvoraIeCOQ/qrjlc36nsl2UQQAg84Ubrrw21795DuXfol/7WJCF8/ynk7aVroB7tyBMAZPhrh
4i6XITef5RdQFCYK+zuyPjBpftpziE9yXqElKt1K2BqYDoCvhtRHA3XM9nLmFtOsaR2KnbK+aE2t
WF1WPRTPs4wKSs683ErQjekpC2Q7oFEMmvMfrKClExofSnCufUEbrinSlXprHAaU4pNe8/UeG1Yu
wNwmWSxlxOJrMFadDXJylTShcjerqX9S5edFXzTo2pt6LV8LB7GxvcJFN8LFFRXre9nntGvGW/wU
W90pq41lsXdmIHySF4wxEt7GqJ/oyqUHBNkmtQCHfutCDoMz/U0kIVMwcumLCfGCkWpC2uLhiFXc
6SkrS7s6uEnrQzMUQSMlu8zJ1Pb26NgEX3oeigPZZc9Mk3jIjnQV5yE2X8hCDFRQHfznAcNaTsc4
iwnLdi8tcYWzNOTZy5fOaE5gbRYVEvacJF6R6UE4dcLRaad5pWLqu3BtZ1aPrVo5jD4sbhK2tli9
WoMdF0v8Dpj2EPzG1lSDggZbQMoZgtVh1ZpscpoURcGgLy9qidc7d7HfT/s3JxJiFkvhmwhGkWBf
XE/1q6vfAqmfSu4NhJ5k/i/d95nO+22xIcHmraMCYFl/0SteNXg5QcvGE0CKKnLwP8d+S0c6+ivB
AbE1YBlpEUDBGLY0C5kN/Kc1B5FwnixEILAH9smwRnAIXxffIVuOHNttRU4KlSsBEVMO4I/rg3my
YqRWukRFQ59bwY7Fjk0WvDd2aLycUESwY9gvBx/SBph9P3Yeg4MstOYrBcj1yAqIli+BL8LtQ6cp
PpSgtunQ/UdTcJgRbxC82OPdx3HY0JnDqJ/j6C39BZWUzQXijOqPJcQ+87m9jVz2ksJdYyBRUww6
rwS6WhABowDYt1pK/V1dY921tthFoOEAb0rSQAgTIaIZIm34rRZR9uKjCCvXcshuHT9mzvX3XJD0
bz8yatAi5kCpRzaXJeWuTbt6bQc18lwMt32TGldYTGVx1ajn8O96C0U+EPrfTx1ra/0bD5p9pPYq
ohudVsCS/Ei8ReKiIw/6HliiI5Nx56tgK1hwy4qjfHs8i4LkK3WRkx7m0F+srIgYsN6zilEVZ9tJ
8mUxactNY0MlOKaJBQBXr29SlxAQeTTuVPOScn19/Yh5IcdDM7oE8V5MEzNgcRRWTWhUv6ucMCa1
unvPhf2LLJ85y+gAv1S5GD5LErtOqZIBxWABwU7kX5LY3tP8ESgzWAG9JQRDfwqs3fwP9oIkcrzE
ufSVdADiTmuLfVrNlNCZJLqYtYLhUt2qHIrsO91IjKLbmDFvcq6HhKGiG/zuY1G7z+1rnJvO00Gf
xBsUOYb8Ny7FC9opC2gQH2w6L/V8rAC8/KIKwX2rEGdxOzRXI276ONlSyC8jz2YApwDP8q0Mj7cW
E0nLnYsIOYsDs93t4FwCewzYWfPLnGjDbFQvjrjD1V8XyT4dGPrJ/Cf4jYtDHhfRJvadJrXlQk0i
svIWOtQc2XkIzibPENoIJEjICkcp5VTJkwSQVxwc+Kji3fubxwmNYMQ970jQWO0nmvYuRqX+9fPN
0sB2EaaH36e7jCMlmcxgwXvIbxEMQyT5jEy3ykufbHOH86H2qLyMI1zd7m61i4S0i55yjfH/zS/x
oOGP77Qq4thIHeI/IT6Mxc+P0UsuS92+BGALRcLc9INMojDvZ2ECHemODMTfOhqwuyQrGr1Z9DEU
Pp7F9aah8L4s+W6jzMnZYOfSTGcW+hNMIg6iXd7fn7GAaFChcKj7liaEGh9SgOUIepRictY/9UGU
wObvCINTeJMRgY+NS45zvmNcFo7p9hlfroghZZX6sjkHFOHXXvmJOM8DyOfhndqC+sRKyMyG71i7
9ZxWuZDMjkUhh2+pPPYng2udRgDgYLNR7b8jAPaHYi9ETaJb7lDjMrcQ6wP4ZblJbVOKEz7ctltO
XeJAav5DceFTUPI6kzeC50Ny53RCUVE38xenUaGLUZsAnrTDLlIa1uH+A0XReJfZ2I2uKr25sms1
JU8RyFHCY6FYkMunKIc2iIAINjnw8vuFADAdKVprfirq4XWudQukpEP0V4YGAmMgwCBruR5cTRhe
BjM9tzKzNbFMyXEOamp9Yv2sgL+HKlViqRZ5viSfhKDeZifb6JjjXgVie8V8R52q7ezToIWrDUb2
LjdKDF+sBFU0yj/llFOENQsP6GdfmTKWU1dH4K+fmX5t4A5Fz8tXrkchqc3tdBlkWCRQ1KooullX
tGNc/oEfi/sy2tt7X3IoSL5POnNRMiDMS2tpa4DbA/xPIqWOTxKVNqv4GRjwFNxpSqQJVBcTeIMR
XMxV3RbxcbhBHsA/ZxXXG5YU+VLuXpEkLQqAG5sgVf1JaIKs2JV+nvsWAJyEDe8wFStAIP7RJHLI
mvly/qyssPW7ZQTuKdLrA+h3jgmWHu2VgAL17iQkmA/LnkVtfTEYiaJi1qa/X+CDRrVTg1y3ud2o
K7tEvIc2+cuQmpTF3t5NT/D4XCyEhNPJlMwVJmbd1SGdAaJnky3i6zygvie1W5dZXlpUL0Z+4WnI
izCA/hPDJxyuIW0aoWJHzYvLM++pxhlJqBfZl1cr4zU4l8MkEbpJJK4b0TK+FjBXDrEdVDwDnkoo
9MuaQN3b3r+9BZ44zy0NGdSdobGdRPne+q1tV94uYeA4PjR+Z+3H6ImsGhgatp8wZloMNSRwWC6v
cOiCjDSR5zAr9p6oGqSceqs+5d4hEFfs1RrFc6rkLM8l0MbZ0fx3mz2/JJcvzFBhgI4HSMlB/+JW
ZmZgkKw7pwwHL/XbXOmr5BnPU7rpj0LKsV4Mh3y+qFy705/sYVofU/PSYPIHdwhTvbEMahsJBQzy
bnW3Y4DrrYR/C5UoPkzn/Eaxbil/8bxuryQNxHyrmhJmZXsEPbiStmjRoUi0vixHMqjH32PVDS36
OMlqkB6AteomSS7e+x91zYJHabfgUnSck5S3B5oOvASSgoPw/04j3Yakdf0jUQjw4KBZ+qgGZFl6
hLDyDuYmIpJ8vPlqasokkZl3jTEnlqyqHbZ6RIYDkjD2HBsIHrDx2FT9xkj6w8/wU5p5kq555g02
NqjhrdM5CV14KxAkU/gi3F6aRPU4L6G5yVbdCBPL3V3nGuQ87w2xfjbzwjh905vOVsFG3hFWaCdU
iq2TyWV+qwrI+bkRhvRIpdUca2Pyiwk1NsPFQ+n/q9+/Ty+y834IT2FfziTJ4MSeUyEqf/8+mDuS
mueyy0gT7dcL3GFzyu5KykKpPa2eGY8xCiq7aB2tP6i+blTqGOaURB2S0chdY5pfS6I77budghXv
49SfZ/2vc5dllvpV72cQAnOo0N3r3aKAJxIP5kIyfoWuCupYsjiuO+bx8eLHXY2kMT4mFtbpN19p
xriuYy03Ija9CRCsw7a3ui1L4yF+/ITxE/VMyYR7bIVXzv3Rone6XNTp00kEXYXO5p4CFF18U5VH
PlB4V1lEFyahgsa4e26BHfhje7bwes0QR3jfROMeby7Do3Q58jYTlqQD8KpkqkeSCdGN3vieEVpU
mDM2DzV/08TV5tn0bJD/q/ijJ59XFpO/ZSa21C8eU3pHOJMNey+vHNsxALiqe4WuiRY+Xr08eLOB
OLaQmUnnrvLut0drY2Ah0ZZ3yyeqwVSYl+jZwf9MFTMpfhAMtg6HvAmtdcRC3BivFxmLJ0imMu5q
kPfrdwdfqlbQt1qVtEF0h+ovgRAWPhsYL2X/vNbB8roqpmxi1tE7sX/WeS0Fp58jD1LZCWwVLFcV
1wpTiyfJpX/ggyCy62Gv9C9E/mfcAd9FaF/REgyIxF49YdUA1Xfo6n5w268QhFKAwHeyiI1exlgJ
T+oxZK96P9ypitXjIqAMt+3W7FhupA+yzog9Jsehar2aRNAOq74xdJVZxaeIfdQRsXT8evVitDBd
pEjocvL1gz+DvyJ9vk2nsH/YFgkr4WbUVWS918bhb68a7KU1dtaEkHkEzOAxRe03zUgZdycky8Hc
aSN4wRwDdLAGye/i5PzJXLh063zeORMb82voKMoTUKJDzZGgIhYDr8AOZ+uWb9KA7pBdnTYJ113Z
6x91A02+3xXKxYatfBFzNJ+BRP8nEtdeI6Nx63Ie3nURAkOCHo0jJqyf+qmS+/EqAU8PFL4CyDmP
WLl0MXU+S0pJODBVPX3WPk7oFGRDryH8CtD2bTE7lSOdEdk5iej2LeR/691lXxuut6ccuoAe0uFz
IN1XszbCeuyRsH4Rgv8W7x5J/EyzlHpZoJ/Wpl7rYUFjoYvkVcVnf5Rat1VhsFfPQHpZ8hAtkcPT
y8EcHSBhojzi8CBsHfc5pODxsMcTRyC7KnP/4XvRuX88TbFSf5u7p3YpWxohdoN/wt17Dqvn9ips
HBihcRMuSlUR4AdyMUxMD+2hdgFPm013MshnWShecZHwwOP7W+fLnK5mo0OhtU6yPwd34TKQpw7w
bNAiL2fEdnck9CXbn0cZSjsytd1s/ViR+9xuOnulVrcibw6B+5i1eD1LLrZMChh3HROHxDaSJ6rK
JTzHuvcc+v5N3AicabFKG0Q8zTQ7J76T5c+oBl3Nst6w8TChn8DGzRRfTaVaVH7etsIoYzNJhrvS
gDpscnww+GkCZAqol+lfDmfVjooY8Q0PyrT0t2D1i1DublpSVMeavjKK0yCBFf6st94QlinV4bH/
Yl6frQbkbE9XysOmHZr3vv7tCYdWQbFiDbASIXGf4LBHoFwWdxXtUkJJHgnQiR0b0IiCmdYQP1yb
pf1oKboaBxPyMqV8fvDXTpRlL+Q0Dymbqp8mS7Y8VvBo7CVGHlQKfkvZEhNETxOgQ+uEiCD5OxLs
K+tR5r9bi0nq8Kng1vsm3xKIqbVynYcwP9qPUGKnu/YH7MZFjxJSDVvDxzmYoUWtr5jWElm74WY7
WmM3zEOikrEHtbsDbjXjqmf0RxlqSB7gZ9PB83IoM1N4dVdYP189058y6ENd1dqWD8XzOMzZGrmf
PtBNwplEn2X6owqP/LsexySATfqlF5MAGrgqW3vIr2+XGSEk+IBFKZLMLvwC+xSW70fcqd4r5NiE
NpZPf/Xbt+iJYVQkWpaITIx6nkcwBqtvFEoM9AYoelApSdQRxb7qu51rRhFAOryjESm4Xzt7+JE1
Un7taS0Hg0ZJyN7T1gFMeEGkf0U4qlntcrVdYP1PaQNe07jVYeARoZqG6pTh4Uq29oqWtzMa5Uh/
7PqGFO/25ykEkp0LlCFbI0HlsIZQTmiPkK+pdlKMNSqLd0unN8wOxNEIdrozmPK7k1BRqmYH2+bz
3BBtXIEv8rXlFmPkWlJfU48xRysa/XwPZH/eO17PLJ/N4KWKUhDX8da+zY4jyZ0CNXbWokiky+KO
AYuQI4/QCVCygLTB7eEnyw4Sh8Y+3BqB7flCyi4zEkaDWJzPq7wA6oV9e1tOEcipi0d3u3TfTveW
CubhS9Fw7JmaIB4lG3xZG2PqUhkCdqFrZdbYSb6DAq1FZ6PJS0xqOxP44gIj2dQkGMNQBz0eOuWh
qzHXR3H8XqX6fsx0Cixmxb4uYntGMV2yR0CliriowAxIqAbA2gtD0BtarGp5dl56sqC+jG3qtm9P
g5SzNAv4aIkeVmIXkQOK3RJb7NhQNn+uCputiA3jQlGPV4nXJcz5sF8ZCCqfDn/i1+C2gWQhjcXg
Z3wsiLdXWVhYWZp8/Og8dWLN5QZpI8DwbW1nh7isLjyrxxf4YRbccICNV4hKG3VRa2IetNij3f8x
n4jlB39/jxNnDBr28xtRdZ66ZD/MSeG0t2hpuu7U8zB1B8WWOEArGV4ViKoQ2C8v9bCnQz+Wd/pr
28bIDAPK3fbrmQs3qDN77+2UEF/aD9yipZFzJ0n8KOKrkoO6vyoJfjnEkOpYn+eAyjjOlAzF7ZS1
jIE6nUowCAPaCvnKG7ySLuvkkXh7un6gPP14M2Gxoz2CGz9giyBGo/iv01PyJUTpEC8Qx48BOIcH
eXGknGQDTsDtw8aKKg+5+8F8aBy0sWfnTTxQF0f2VQfA06al2cEy3NC3G4Rx1m7Glmc0YBMmlc5b
a91eyAIW79sVbV/8a6W3bg2agU1K/IZzuBBorQAY+HmbHMfNWJvdQa0/AprQ0t3WN+FePkcKrIga
ezjUFG/kxyk/19wLk/tS2q15I3Fsc3lxZMTXERN/ywD9CPvM+DbYgyKOipakmHV6UMRR2Ey0kv/t
c//XhIQQpMK+3cPrwmPIgQ6VNGYR7Gkd9d1++9f5V88YY34VmVKXh+wciEsEPl9pXgznTK/LASvF
LjIuwJ3oAv97nsXv6b4hGm7bQ1kd/gN9W1ADaLkcp47Cd0BAiv4Gbxj1ZzM+U1LNKc+qb7ZECFzF
MkX5UIUqW78KDtU7lb9QPnfAzYl3eHCzmXFb+BuXIiNjaAHgcbJmxu2t6k9dtU2girrLw+s3YyeN
9mPLprn09+AEoU5r0KvEC71s1ed+F/3IZYAMNzvn/DJCB4mjnDROAS02+0xTfwwVBjVOQVPtPMzG
GG4tZyHhPRlxLOPjHAKrOLCqBihcCT0Ogebo/uhKtpbzMvzSPLplZABaqqAUDVIhpjDROL6U06Ah
nSNdcSUo10GHIWE9jtQLI/o6ONZKMF34iMB9/9pIqbA5ehDfti/RUoZoINM1vlDXhtuqOPb09no3
UFoXSM+UDCDHS9+4lxaZiUOfhl9TzHj25qKOn3jhJv/gzDC5ye5A79pYcnnCN+mlLUKrxjLiVSLh
gauH1FXxaq056R5sjrtm7JvDnU4LhZ0+VRJwq0129MKu5PWFt69iSupW0x5dKUdFYB8TMrj+lqIF
+xhpO29mSVn9+RsO3O3RSavcjMxoHwaVvxN1ko0R5B0I5QzBqzdswHq2mC17or23PxDblWtJtRmG
x6a8JSZoXWBPGn35GQbrvpGkfm+VF7AcEYnUqTi8Wn+2M3LwSegfgYCd10goJza6bOlHuOWsE0Kb
mEcDms9IIkStqGn+yu27MwQf/8ozX/x+V043LH3EnKO+n32l3aammxfh294tnWaLNZI0fskirRwH
wNCz+SHjVahT9RGAbP3/HuFNPrci6KJoetCxJ4hhHDJ6v0F7Jp4EWGTfTH6Xl1HyJrJ8BvKfkNOC
hM3BuK4MPdZxSI8aFEccJl8dGs71t6JuQwSbF6/lUoTvv1h/IgATAcvJ9NsNUAJolP/w8nwZuEQ6
m7TAF5UcMGklHozwp93r7UTIeMF1RFgQ9SR+VsaMb9HItFo4jtJkjKb+dgVQHSDLlvy/eGM9lsGD
6BeO9S78R10KStFLKIOZC2S04JUV3UcHMMPtRHM6I2N+eby0ijs6JtuKYsohI3Ebse2lIUzqQw3c
CpMNqn1UZ20MEbb5OoCctGMmnd9A9H36b1nCHp9UBcPyzha2CRNtaXstWhm2hMZBN5Xzk4DL3x3a
lNgqxQlJt2Q0272WKVHbyXt5OgZH+I3r+Wb7uxXRrl6sBv+S4TesuE+vujKYVl0YfAqsqcLJmTLc
vTCdSgssp5+Z8pJGZFDocW3GfvlinBx91tClYXk+cRtSrUA5QNWjj6fRuNSO2x4hDVxSayGEy/Xk
EHP89+spWeYYWD5N+uiIdwPlG8pn6sW2E42/9vBBt39kMRP8eoaI+I+EB1uvHZPVBH1qdlO3kGhZ
TBdI/0NVk+ZxNUBAuUtrjnUpaoo+LeGIqxxBvhT6/PRMsVD5LwlqqSGwFCL7W/OjW4NUhb6b13EU
Exm/iyAFt9tp/u2tW+PKktM1g1/T4/WI5qXx3U+XA2gugT/Y8pCYPS1UIef9bfesPA0d9Gdwc9PR
kapi2QVFN03jLGvTo2E+jZ5p6Z4AqqO5rWUaNgF55D1Hsu7g+cu2Q7tKEALMH4oyVoj/b+yoOTTa
IDj/AzMoRNBmHZLUB6tk1jGmoWMaxSMFEZL50c+OZs8K7g0QZjvBpgtGKfJeZ333TWi8XtZdDkqJ
UNU8ibJgJMg3xbXwgFIECwUb362H+MeG7T/miQ6EQWVrAAD8P5m9ztCawfUYmJ+Zj4EfpqojwEGM
UdjVkZCko1K/gKA2YBPlocHL7htIBCfue1ZKSaQ/csMHr4+Ix31JppIShhbOFTHKKRdwdD3Q2Xe6
U0UGUma0BM+5hdvI+fct7AWQRgv5h1iXoPlptE9xYv1hvXJLf1EEfPb0WozpY2jyDDNxQVIimKGJ
MP8zn/KeQ+rxaHIENXm5ieoB5X6nWWxIHTwwvaxRxaJewW3qrvuvq5ofeysQHTWtFItwKj/AO10k
fKeRI1VEz4SGUcohsKTSOOiEKIUOLM3365y8efEea+MvtzDIg5vgtUEpa3kQud+Devdgv7d99QbM
MfO6ewUWK48cueZeqrBkhXqArxbHAMwR8pdpqHkbKT8WRS/IsQVv2uPKgluu0z7mlfwDIrvbbcXG
1RA5E1YxBnMYbo/jqrDwkxE+JZ8tfkhHJMb/ixhSphjm73pK5caFg1UWMow9PLAXSLJlvTJSRBnH
xLOg9H0+BObg9Vm2LSTHIlpHyX3gZvgrTuJACL014tHpk2/lr6XlhAuIwVcCkaZfvEOwAqmkkaqK
piZ3sms8EFYu8UugOkSnfawYlnBnxD4ivF4cg18a9/z0aRr8cMmcIZzAu2gF9EKjjkngcxy53alG
jrmnmqp3I3Z61frnoM4stIdh4gR3jZWDhqOr96gEDrA+3sFP1a9R6Seq3OKkJ7t6A6dHzq6oQFNt
642yY7dMDwfcdDdTeaDISL58oco3mjubgCfnX7nbBs0SOsPuuT6tRCr1T9EJPWkuyHbLCmEMwuIs
hhbjNDoLMBQQrh2PKr58BHS0apc3b8FPAvgFxZe+8TV405LhslJUK3om/Bp436zfKRdLQXfhdEXN
2ReDEZktKuQjJw5ZWbkh2zBySGOTb1Cs5u+hBl0owXLpiKhimfAN12Dc26zD6YGjlg6TkXKGxoTH
HhXjV3F2rqugC2T/D/ZM2TdTDnTm8OUfqZNgxMRChLQZKc3UBwlkFiHZg4oFpbf7t54yCYvvzqPb
1o5P+YRuVDqdgTdnCRIxzV0aODgtQNiZKbe7v6G6dj8uS5SCxDLFTNEEFxCc3D6CUqvFQyy/MInm
xYuucThq964Jv0ziGZG9pDlCK+EEMDBb8Z6I6KUsGcdU7q+9WeGDahxicKeWxNZDIfAFJL01Ahxs
1e//RkEwityU4ZsO4me4JRDfCb1CAodcGjewheShYeBKd8Ly0GyNfq5k5qgPgfULaqAiqDloYOhY
TzT3watFgNhxD6AxlF+ck0ioCHpiZ23ObBAFbmAy/am8+CoqE+FXelSFTTdB8SwMZ4e7J+TjEJdH
KUKDrj694ecDV9nU+dK2ku/oIwwC/NKkOtVT7Brca8hh2PDbcJ2sdb8EezLTYZCZ7FxRXiemEh2V
sg7yTA5RsQj4PCtYuwuA/Q4ZdLuYYJzm84g7DXgMAtQpjWQq29gZrtJeqhkkihSVK/04LfWRt5/E
yomOjI6D5+y6relhqxieOWQtV/F5yw2rOPAF9sgQsF7IA3Y9sYodXpoXRrRic2A/GVWxWtjnZiTQ
rWvnTHQdyXx9fXKhIXf0XY9QUmUt2ypOLhdRlEpAoc90AYzaHqiSzB/XsSvsmjq2Nj67EO6w84/v
Nv3/Kv7eblZN9mOZLHhwE8FoJpoFMnZJCV1xcMEHrs39gwj0mu1zpYzLq79vc4GBETNkEPb23DU8
LRIHvP6wcfsfDfBa7ao+SzXCszm8ZNZyh9IEJhmEdQB46Jt6lnQj9RrBmBX9AtmNPLxapj+ms1Ku
x/LL+MHClPxInv4k4esRzM+75JEku9UOFPa6VIC6+Lp6TsGyTzNB6YQ+OskZjrOzQddWi3b7VtZr
m7fZeBIbsqGP3V1Xz6qMTN91Bde7LssD4dLBP0VXQzKi5ASAIcg+cY9kBhBmZkFTPVTErIBJ0Ty2
GY2ylSL3TuyV7FPoUC880AeCgScFk+mKZTypeQ6PRaj+NWNcdF5Sm2g7ZWuh0q9bo4khYKZXogsH
VlVi1P7qZW3FBLXaHooizdcffWUh9XocrS84sKVMtLYrsDTxpfNlmy5yzjKEFRBCT6yefq8iVeRB
PPhq+SIE4dfd7W+pWlJEipirJ1wsF6eebCu8YefWr/Ce/kTC/V99xx/YrFFEltEpCdRgggw7tNv2
gkDuu0uwpbnBil8ZbAEhF8WNxlu0j200jEFG9NvD+tVTluW02ZFYyOn3S2ca9l2J2FfB0R5Zk1Yz
HdcKpdCM3jh6gH6ZFdn8qv8rR1vCawp8hvdu9yDZ+6b6U4M1NMzIkDe9xQlOqH595gstGJjjfPVZ
+3uiBg9wSZOSMHGDMQc80b9hpwGh7eQBn3PTmeo6b3WeI+GRAwhymC3mGONMLhmHRYVS57IBPe6N
WyWsB0wDZLz7Pw7Md5Uez0ODfqpte2H9MeSKsG9huWl2MhsFbsqflk6oMbnOV9im15dICq2lliHU
kMaJKlQv9QFVqpeCXTkbn/SrQfzOmv3MWpI6pi+s+QOw/uHBj4l28ZROH0F/oLYWmy5q8BBOHh2o
Qjvs1/0qtj7ZOfpJa1ThtKfj+dLkzWgRS/xY5I+fcUqFLQYMVJXp7p5wuafcnVKo9DkC4JB6WZdz
7rRFWO/CQjRuKLKFyqLR/JfxnuRghyGKjT87WSoeLbbWEagoyfWMX358mSQ98GffUQYuIO1v2dtH
OdSxwC+AToj6E+Z66kkeBfUqSvzsfxWetD4VHFwgnaAbI5mXdYB0VP/xDR7K5IFtWfw3ItJsAcYV
sLiin7TcojN9S6L4ZNuXSblSxYbbSFGGXxri18nVcesspi+Y7o6aD50fe6iTOEJM/9B5DqUiv/La
sZQGoRbhq7hcVh3ivHBhNTfHNvrm8Y3PztifA3MarSVAPUVPaEcjwysbOToSlsX0eBZKywhFpi9R
w7xDIiY/h9lfNGdSgr/1+W1GjIrVNLJio5XcOkPtVFGB+wSn7+jUdQADbqtCSc6pdfT1fxyFb8zZ
GCfQjk0NGsLigUmnwi4kM8RCKnDx/LESxq1PngvpJdgAwo8fd03nnX2rDbBvJx50/PKvcEKszAug
OVrDiphuqnheWFPiGhas2PAjlHGwNZTSg4/kaxdzVD84ndtmetbCXRAw2RR0ZLj/f8s3ht5XdEF4
CT10CpDy+IGrnczC9Oig1U/phRm/G/QnfWYiSaPNHW6E3rtMKIvw4754Irk9J8LwLiQ44BBeUNwn
PCxkfW656SNI75mY3rDed90Lr/dTTh2VtLbRrZRt9bL/BUfe5Hrt9seBsc1qmSiPO97dCa7r+su6
6RvloD1VefumjMxxgg74LzpRHw2JbDeyZxXMUP8kK3JsZnSHXbPF/ybNUA/jQyWbJV6UG9yqWDuU
MjidMJEvXLkTtt0kIaYJsv1/YvggCKWd8sW/HfcPX4rLkCsr0DjaEufuNGwEXlBG+kU8RpLdTY4v
bylai7pPbFjLoolTKRPx0Asw+zPh9RTcy5F0OJcaKqZM05CmcNKRptNsM9cxe5ud59KTgIq6e+tz
DyVe6xyegdwsyr/eK0gXXhdmy/ToEd3i7JV3hZnVx6WfZx/MmQCyQOU9+lB9/Oo+8x1gnD1mM3A4
81etf5CMgzR3rSHkXAtQJHfteLnRwSysBrK2JIKxcVzoGjaILJZQZhDw60j9eTLgXRjT5AwcBrnR
U8mdtd/NZyzgYbFplsMhQ8N6UPldezYKol/VZSAL2SV3xIFX+8Flr6Rkb4UFOARUQCyYy2z39IWX
+1U+ED6TPfrSb9h+a+UqCtchOO7D7Ry79gKiZ7HsUbpGYMmkkkFRfwfPmPmjFWBIvmRuHoDYhuFJ
/7t+JkU8FTJISrHGOorvgLjlK5Zy1Oa+coNdLQpmtMX4qQCXQw1M82dhCcELq3B4iPNTzybM8dqb
RPCJMEAvVGfVdTPJZI+w7Htr8YWA0TYqbTeoQoB2dRlj8f3qnd4aawNc3bEXvB4pugVET0hZTTxr
FPCkKbkGus8FBpesd6m1CHbHACX0m9X7vHVgHyHfJQEfr+1GuggaL4/aIpYjdfJCwD2vlGVnXFHc
IkNZ1qtuKierdLotYpQJQ5l4Xp3MdJ4O6WsjTpHjbDzbXeuGCBars21hrQjlTYScGBLKglvunyWh
kgmdYC7hmmhndndV0XffQhe3LRcmFRjXlFPj51M+a5Aq1YOldCP59rJhdRoavjuW8AhdA3Th0ZvQ
oiHzTzea/qq1ppbcPw65BEz6Q3A2P0kCQGy1/U501ZOqA99hTsV4o2K2aEtJHmFgZD8NDWHFmyYm
JJW0ht5L3UXLXPLAxKsIjao3Yh9kr2YMNwHa32fL0CK8Rp6JJCV/g2WxUsHWcNPIlBSCx/pNmQ4x
UGFBG02HJLavXi0TxS9wfrTjXM3G/DvGpq4Qyq/S0fV1zx9eaK8YuI7MX5yObN64aGO+bDXrfpxY
baOE3kWaGbHFdBu1RscnFsydGKwZCgScgNn1y3/6s5ipqW1xpyohq/FoQQuQQgP4A0AXgosLq955
nEo0eJulRp719VkN1DmYdtvbFNqFHqXTl1LG0qWkgEtG0+/r/J6blhMAYGtohQui7Qqpc2W0CXSn
xsTT4YYMbrfgRWhqaEh7ihO6mlO6QqsP0pzwL0kjBeVLWw5SBmc2RULGVwE632IRati72b7BkL8p
heD5YQZs2ehGSQDfw7PaMUbOlt+qsCHHHfI83ndOtSlTcxd1VednYO1YlRBOQ5AU2Z1TLt8amEcr
joDEdCxAM3lQVM6e495vMNpPykGU3E6rFmuDugytqN42b67FMBDKqISDrAbSQWu1WqK6OyOck0Ug
2jfTUgskLwAUQLbatXraY+qfWvfGf7njoZUniFSMGtGJce7NEWupu2rVqpMqOvgCMCA1zcAjZWMT
qVS5hlKAuIxXJwWK0btJIP4UtUVMiPiIbluHoozeLXLNSTdU8DFih/kr72G/xGti0CglIa6UwDoV
0ulPUxp1O+nVMX7bGe41fa86myu8w1hDNVRKkUTEALeBhXvN7dJUd1WcO8cT/eL4Wo3b+XKZgugt
Kh4jF/TC/oNFoZkT57mIi+7MMRyy2fNuIfBbS/QoJRf2Q0taEodwuO44EzLFrVFrNGk+9R2RPN0A
dBNjhJpLAwHfwtXxzrJNsbZLu3iUco8Ouog9QoXsaiPbHrQPgFfPsCRyz/EIB3gGrN7pVN2UJEt0
sWAUj2xqeYraNEPHunDucXNawRwUZCAFhd0SMRideWSnYew/WmgO8d/ls8TEKfLDZUy1bnma1kNd
Xp/SVnUrCPDGiQBGCfI4Wh6gNnLV6xCjnvEymTbc+LXn+A6K7WDaZxalfkjkz0vVcAXbEGjIP7E2
yTVEqpF1qNS0qx63j2c6FXr7UNUQTGGdr3L1aA6O809MLLwWnprTFostt493hXKNU8KJCpV5JWDZ
9gzpOBfEtMv1gYyPZCN27SpgdlhRZrzOPZdDnvwbQiTgYZRYMYGgDYem7X8MmUPcQqFuVLD7QtkX
CITse9Vj7Aip5RvQabBpDbHYGsyV38rPx/nEU3iHSSJrSsN5d9OsCoKQib5ILbOTZuUlhXON+i9T
BbQIxWUt3jQrlW+B45krbs2h6XAasjRvWWfdNITG9NMl57moWshD2ZLEgMmhffy2eSDFZFlgwJv1
p3pOyLGyuCRe0BbeouFA0fKRCd44ano4oO+6j26AxSTgM4gBo1kMCs9TlCFEXfuFiboiQMzjoImU
4vOMOaQ1H0lTNMVW1vKVEtkbPddVtxdWikVFZEGLScbh96ZUSjAPtkYoLMEopWGsV9LdErOS2U7u
fo0Bmg2cS8mZYizfkn6VUCKZE2761loYVIgVW+K4mwP39h4VBCA5bSIMBpMJeGgmL+6wHJFGvT6U
5LoFwWbB3CSwAYFWmiZzTl/WHGyt0PRdaqEKL+dS9BoN5CyBptJQEbrEJuqjupa1+e/8kEomLtuW
aiigvrhMJ5AdiRPAzIuaqCoG52HQcpBRJeECIlwv95u2KkNHmhTYEGqHgfP+hk4A6Px+1SOpms0t
LzDwKpqP9IeYsFOM3CosW42nD0A8AvkqLcMJ0T5dYPJVfukcIh8C34f2rT6piu1AQEhedkMYBxXP
6haBrpmNAqZGEXWs9mxCeq21bjndX38QxA2dOxy07NzU1Y5GuV8dUgqaqqd33Li2etl1kWUxHXjA
A2rvxLEuWla6kKXaCyUULht+bJ2eF/nYufXHW4opoGyuY1F3oa7++AHHvA1U7VTWvlB1EluC75eh
0wfmpyjtX52FP37RJq6R5BLbCKomQ9KCUe9O4WnISfPpBWUcaiBOmMSpJ9tduB8KxbEqmzmuUatP
rozK1uBITAWo9jEAgpqM/JDxkFO0qR3iRyHG3Dp+FSvP4yHvApt3IM6+Y6sSsLfdGwLI2mR5Wm46
4+v8WwG5WUFur+z4bHRqvl/N6D1gWSkQhDHcsIMk6gNTRSmkvacy60i7fhR6iCRZ7B7Il7ZOJPbL
YYKWqr9R3WVB1lkrFY+xotABuC76R/FZbxDpfaoKPJyLNFEL9pQRfJrpZ9xCc1l2cZp7ghxa30mc
qZ8aam9UwUYZEDKrbydvC1Nxlvarr2owURwdz7G/UE2fro/ncQAVYKATZxkaOA1iTYQn2jHk2nG2
h46pL2n0y1IpF9nRCacIy82G0hDUAFjiTrFNxb5DQ4ZwWWsN5P3fZgOiHiDOhO125xU4VNk5dkHZ
AMOU1t4wIju+tFHD3G/b6Mao64EDGHwkdx1wmLAdaJ6x0JyoDS6QDu8GADTeKl/tO9gCaxUX7bev
Hj/PcUy4LsnY62CrsxNGQWEjsXPBIsSta4EeN47EyjJvFvT/cnK+ZWp4cfMj65Nm22okosYySCyz
USoNzgXmrM0oTDacKWkRJvFvtwcycaMYjJ+jsqQsOXwiRVv9rqTPE8GmJKWhjVqg/vu2AYC1vXAj
yXWmsC/xal5Cb5MVqFg7EiFY2yIuSqLU09mZQU46joq33ppu2L5wZLxUyPjpCYj8qjpBH0vk3OAD
iWTDCLJKCn/ip0Y4ownSJJRz/KSd5T+qtPwXHiCgjCcTlmtsC3zQZ1tEHRUUysmS0B2paQz/hOU2
848+PT7Cua9okGhi8+rRhswK2Cv1jzY1qbTj+Y1j3UclGXYOXcRYstoBDC8WIzL/e5lo17LdXw1o
fEZ5MGvQgZfc/BOYbnVWHICRb4XC5wqL6dq/yJ7n9GVNVezw7dC2uz9YKK2DrYuJtkdHkDW/sOcS
pXkhS+6ybKpIxuAsT/vXQWQNzaVHCkOYJMy8ZCgGsBaFo0lqkABvg/tFQFvZSByVWEgWoHkU7JHL
VXOR6GNwulprF5i6Dc2ha6pNwRofjajTXSo9HYRSz6vFBJjRellTVcD1egoRVqpv2dQ5/2F8tvwJ
t0L/7TGXL2cBxNhQxhD7x1RsZ+Z+0bzJbEFCitH4uCK7dWDX03liXAJnkDKKrAAKEhAQqD/YVwKG
PeD/1dwdQLwjvq1eX54gGN25QtMLf3EYeH60x68Necmamb6rpQVUDLJnExK1GDsnCYUQQZ1lyvPv
Km5pOXIr6KdYb7ZfJXG9pd2vpXvAkeoehUNm8tVRKmibWIMJjSVw49cvtf8uS2/wdO1ZbByoloeP
LAf2b00j5BEq6YdSg+faPpl6SpDjAwj4Ci60gW+SQ6zjogPnuicAR0HRiSgemgQKrJ8bMPyuYkVR
HiIbF+kJGjh/cyQ7ZwnPr3zslADB3NYmUJscLqZx2mCIZfoFYo/TdmW8/kCcFGypYQSjhGKE6WU6
DfSiLMFZhiog9M69oTLvWQcRNXeJ6GChnmNQAFKluU3QVEI4JltPHMfk1k79ysXO2d5ULfXHC/U5
1DQ6eeIaUNd3UMF1sKh6xp4m6LDJCS89SsLssOUtiUBZ62AU9WaqDdkkrZNoVb/JrtsC7Gc/b7Ji
Dr2YozlmPtO9OfnZ4DAeTwjbKLqgKLJhoqvZYDkdyz5M0U6ag8SuPXOMBqu3DUvqF6HTtRQDpgJn
fAizaSZvuQYXmC4Wyl5rlacFjh2aEm4unr1P9b0mRSZgnkymVhSmj6kTr/i8aEsrI9MxZoS/wnnm
U5LkdXAqnnRQPvdHqyti5aLeTl3unn0mQgbGv93YkwDQD2iXMoML20JIEdDS9k0DWVJZ4m7esF/l
3H5P3FQvuSrqRKbnzDHaOMmXhF8rM7+DjM5ta3XRYUtxcJFxlpWSfEa/Msht0XqpJHKx635j3HuM
Rd2rYD0LdszL3w8TB6R+Rzv/1DsNeKBk2HNhTuT7epjVpOD7fRF0pITnaWMWAGGEPomVNgjO4+V4
AafvB8048X/7XsST/kK7NZz1H+fu+z5zKR/Q1RSdzdyEIOCAh7tsmfyiFma6eVEPM7+Insbm4SwZ
prftLRt1WfoU5ttImcU3io+QSgMARotUoMuJsffPJIE01JIYsOGPKpHjpFlszOBjztJcqxWaH8sw
UMzQtf2AtgJUJQhLl5U17ynxviTgJhYeZ6rHkPI6FjWhah4v/BSjgGqX2BKcCm/zXsfaezCG86R9
tGPxckAtGFEzNJFrOIO4r46UlrRjuuKKFImH3L0qgsRMwCfi1ZHveAYUstcYC5JD8l5M0FoH4nCT
jlJpaGVpP1FcfsIZUMQEhEQvO5l7/S0hQwD35XiuMCTMmNK0XUISLTlH9OWaWqH/zsBxNVrRTDoI
C3YKRHPghvLvdddiyrz0RoQAELxuPC1wgy627HBt33MImKLnHc7ECYQI8YWhR5IrXahWEaMOmG+b
bTjUJhz35U6F+NPN3BhgOMHMpbL2T3ByESlx6cO1DAIp7KWb9kBmCNlXq35xAQ/+Tmolly5WbjPp
Jhs2kJSLgoN8CY1ZF/dqlgufMiuo5KFkfv8+zTS+KkpTq5YzADtloAPEDN5tqVv93FUAqvpz+ybQ
ql8Ewr61ySSOJUWe2MyOg9WGSofLM84utUorvGNB1S04UhTXXbRTHBodSzr7jZI96VkphvNjq1Jb
5XzLR9lG1xM7HIRQ9M9BsJe15qhGa2z1tFwmgXp0hxH2vO0LVJ/WPLoz1K51qVsiE023QKyoO9gh
vq6CUCyPDuFMbGe/ISzRBfsXFj7u3HTtgqqkl54DtALAko615I61V0Cmo1Amb72YoytlVowtDc6A
sxra/qRKAMy24Nvf2PmwK+6vpb7kMNrIYptEVJEQwBbfP+KOkG+2FgOk85lp337OkAqGpJ2UbJ2a
z6qeQGQHpfOhiiFJvU8Ggh+y353AOtgjsbfoMR1t6ThmTfWSWkj9JLNzPLRpofowK4k3v8tJwh1g
k8iLQUmjc4aTdU53bInA1WNhQXOg64MnocDaW+y5iwMrwWgc8KncJ2vgSFh71T4EfcAah+8Acwen
beyAcnq3+/pNdA05wwcFiyLt2Fb198ayjCfD5BU7g7+gBaLlnOPdi9bCPh2WLtdRCcqXOSdDl4/2
YKnMQABUzqOYwFbm+6mBDl6ADKfTIkn2oyVbGjbiZFvjtOhDHgY7XU5qYoYV0S1YACGL9VoXvjDz
jvpnXA/9dRQ2beYAp/P7BeGZz0i2fUIZWwrmBZyJqtDlDf0k9Y4zIOG+QaiyI/Ehk9g0btWEyIfG
HyZxm9xMLEfxFijNsiFQbUyk+ZVqXY/Nj9nlhFcaBQxby967ojRXLcZH1gFRzO8HA4VAXHCRCQko
PekBrD+um4J77332/1qdGTmi0RBPg74qN8litLykIXnZZGdDG0tdlVqyf6pAbV8/+o0knB0EhN/g
X20R3aJu7QFRml0m+nZwv23Z8BvUqB/5R9CaEfX6XHxvaCvWeUEfI3hhsRBm15SDGLzV5JduPZPm
Z/hpAlcmdgbp73R2MZ35sEp53k1lFuee2dPsvwWfPi0CeqeuYuGTFayEOX5AUPmihyaC26+WnVHa
eTcaAaJGpQN6WgkfdesOanaBfKoWlR2YZDDi6cYtzPU8TWybY+IXgLXBfPgqAUI14qI0V9Iw79Zh
u5Rpp+O9dgoMCLiNGjFPrMCk0kVyzzR4CZ3gzd8YLHk8UdnF19BIMU4Qu5qmMGUS6YLzslukoi7D
tOfezJqXv0EXV5yqVZlA/BJGnCFwB6H0kBGFsmhcW1kt2uLDtGPb608yqyIpjhMz8bzbcsJiRpZh
bNvzdTuptHz5PhNN2T+ZGo6hU9CPiJkW/0xjqhVPWOTvZusNmudIAbIHPAMxTdJemcTQ+SdxtMq8
WnigjujojML5VI41QSjs2Fzw4hagjdCJkphdPTGcDtu9UWQKQjQr/G+Mx6I9m5Awn0NWdTU4kisn
z/qnh6eTyaThygyjup2WkBrAA8iVSgk8xbeneDgEb7T9GEp+OEAtesybT5Q3ndfNmW1X+26InZbm
U7S6SZsdQav+3IamRrDCTFT2fHHMu8Oiydc7zZF0jK+/3T40cKh4IrLcJlNVM8DiK5ZneqdkMQP6
Xa0yqVHwpW+fhwA2bghkD5KukTSCJhjns6FA8SoJpuJhqOMMKv32UpLAgZ+KWzPpFEbsbpImfPib
dHwBBUY6659DVc431i2ez34gMqcKOF/EqdOy/n4R/y5+xz31Rj+YckPPfDRYteXgi3nQIOFH7VgJ
iCp1Xk8gAlOiKi5lgSRdWDSoCh4IKqtrLpPDKfI+5izO4c0H7bQNNeb1YoNWoCxo15pPqlU+tpmM
t1d/GtU3pEPF8lmnbotHBbAOLpQ2ZtjBcYA6Rk6a5g8DL3FkHFNhjVVkCJCBwLZENZIOLR4KIoH7
+Fx4OzaURMQojjyZDvaD6SsI4KcWUdrJavkdf79yS1Ci3HhKZi7NRb0FGpAZomvHeL1UYaLFC3wh
4X3MD5aaf2wbdRbTZHDuOzCbLL2O2GgpVWxzyUuTKEsT22qG8bwM3ojbPkCqxYOrH7BuSf4R5JBU
5n+ZHny2TcOlCQNuAHV1fXyElxHmF8SV43DFcvi+swqnc9l8cfN9cpN3nVxgDgmxIKzvZvyGEg/4
T17IUXWFGt/+Gl6Ks6W1wRiOcZA9Law/nzblH42GgTrD6PKgO1U+ibFkN6u7aMrChS71ksPtTQJT
+6toot1TgRxkiTTVDS8K2uXzmIMUKj4M+sfWKHT17HVt4CXQjOboGFG3Y4++M5MNvVbHZ7wr3hUY
d1dkQxZ4om/UXxez+gsvKAJ1VQ6J3We4GycOM61G5tCRef+OM0cfhVd+aZtNJSD/afdLF4QFd+hJ
k8qmAkBx3vbsGRrwGvE4kQtq7ZVsNdIHgFI0bA37gAj7zzF178dY0J2zLnRJVtATYIxYcjUEYVy9
16cyrCkiFgtsFxwUtdZ3ipVwqikzFsXMA6ufEqdonWsMwjrjQ9xg7ARezkRfF04Ih57cvhQRTHsv
cn5r8gvkjAN8Yq6/t9ZopXHA8brDUU/lmwUBow2FbDq7jcr3DUQ18bCEF+ZB+BGhGbwBvC3ssf0F
OfKagz5rDbJ6OM/X8SW7ZK8zYn1DqrMQ2qZGjeUo6JH6SSPQU0mWI8uZYEEFpXgZaz6rMuV0BjCe
I9/Alg69S4vmTGs0FY+xnHcKWhNhBjFV+O/O9hnXaPm6HnjrCUq7NRWPn4dY3rU3aHe5W20CkOa/
+jn4askoyJ3SF1qPGgydK7iXzO30UmvGdHYsLprtAD4622sXGBTQ6IEsxnlCnI4jjv1UeiDaWR/f
fCxEwKp8zEzgF6rrgs5gSHPg/fbozbxyaPzwbN/6MX9LsKLEbo2VhujhTzlNpyCuoQhzyDmn+DoQ
3Fara07L2wX+RgsxR9o9wlcTYiTctkXPaGc0u8pWd8kx2giW6dZ++mn4/jXGFcDmiDEpVd9DqbDf
xz4Su1xlFYdxtm6HTYcYS/+8XAILwx845DY3KD40dTexuzwuYg0vinHyj+/wcJvrZ1zluDggAZBl
lfrzanbJKVZWIjP6NrR/G3/YU4OZ3uLyWaDkZCnfnsqWKs9RN+RpTMM3mnug5I+Q28DQpTHc7xDv
l2jIR8FcoXnbSuoB4wXh8gLmbZ37vZy4vOJpT9zyftUQ5LLMEYfCIHa/lRc8uZiU/y8Iwi0lPrxN
wJnKW4YPQpuNicyAKlmiUVnCdY7hke3XhC/j16GU9/1D9EjWjkYKmNIQN7+krETCv/5R/pvww50N
JA1pMEXsrs023lLivLxauOZO06a0ITbJ77qZ4Ii0SFERGE3tR+QKM2XPIYbHhboLF2n+4oOcFM15
aotYCPNJf53OLBRNMxdC/kAkIfkaMMuOLJQWTjX47tXi1pGB8GT8RWKLZlAWvRRpN1Y2Zh0MVbaW
jSEx0OIP2aM4ldplTYWR9TztWV7j0kTStZppkVClp9R8vEOL2iV4gGnYuGZuh3gMsiBO6F84JWH7
adBNm0e8j1NTubrMNqhRoo9LKloGbgJeL0hfsywMhFYD5p8BItNzDBKvDM9nc9M7BZ9x2aZSq+9r
B6/IZASNJQMHXLsHV2+atVA2z1Q9EQFx+f9mksIPgrNTYOxs1BpbJJsySNtQc1XwQsTp6HajgsQ/
ec7PU8DW1VjkwYcwkFmMv7TmXiPpz6mLz/L3hfLzf2jxK5FMLwYMrDvzRaDxN3azb+6uAGGf4ZHb
R9zgH2wa5XY+AC2YhFHEGJYByA4pdigzDlCF5BsJUPTajLA7x34Tb3iVig493vbobLqKmhKPLjLg
ggD5n85HTdAGsjK9v3FIaDSOWLfdZ0AlBW58OfGbx29LjpZP2jauRuJLobzz2nblMZl/Tp17fVnW
iTSAFEZnIhHTh340y0fHkdYixYzPj9q0Ne5vqoUuhfosRpjQ5xGfq+S1YR2xeHbRjgVhv4MBqU5c
vomPesyfe9KX/5yXmtdY2uLROTFuaJynz6JGNjpk5oF7+jWiwJNGAzBdSQE02NbbDPYUSlaq54nU
QhL9HWKt9hgEiSNsllDTOT71hbqd1RA3Ctn7b7DqoII6+D2xd9toCKFYiu0EkI+9k8KulYkjMZ37
A6PTlQg6WNZCxUZnn8usFnY0TX8qWE1zCI4MPb2m0ICPusTLMoz/BA9R8Rky4G5Nk/NDW2ocQd7T
yoE5znEDPfAbd4MQEbkzXqEZIiVrS7Uc2b20GnGVFsRoNQj0qVLHmq6xfAGhEp0IiKkgtbznsigk
2y2ZbM8qJ5sNQlbITpE8XQiY2w7b08LqCqItQpgzYvM/1vwAXQd3Nx9mBCl/qQM5oWdLm6cZ+7NE
V1VuvWoZckiz9f8Uvp0YRd9zlb0QIefTfoHscQ93OiEwihHphYws/Dv63tNeEF6MXVF+dcafMSQa
h3EKIZgrIrHX7Gp0Vy8QIQ5SbYOQXcK2TZnpSTKAaV71PD6wS9R5TvNwTlMNlm9vNqa3Crwfpx34
CF6CQzbxCDdUsFqN08zG7DiGmlH1zvSRgYZLag2EXU2nuDQ8t9ZopBRzlXn/BSQSUn2odJ1BZI9l
EMc8aR0FxOBcN2tUA4OPLaqREb6CGlEeNFx6HfsYy3kkqmYv5OTzY0TwtgiJOd6J9FVYmpvncmAN
oHc+y7010RaViZ0iCd2y/Pvl2NYaqRt+i1N8Sfpah08TCOp78Xm0QdYcIz+s9WroE/m2ztIX2RVG
nGOJlZueoPgz34c8lEyqT5Hf7ltTjy1IhDGM/3UdHKAJn3n7886XTaF9K9F6gvc5dYZ8SoQKXbxf
QdcKiEUSgMIP5n3N/JP484Y5bCawj3JPfuVMQn3sqy5mV8lSMmRNPfpAFd37z5EhJC2Zj9IlbEfq
mp0e6GaPquYiB/rXCmMQj6nfei+/DL7QWq3U8rUn7+ChlPYoey0KhjGHkMd9Td6INQshDphNCbSS
QoP1/4R53iHRs3g3hkcyv6HngMXW5JOZVyAJbTq/LcGSmZxYQWGAg6WWgghm2J+MFPhifXY8AOM9
4VFDwYKyy4qg3ZI/kI2MByitymMtQZq+hoipquha6X+0fj6fAR7+DFgTLAww8W/U+Fd1ZOMVeZl6
2QqGDu/onO9GW/jrm4ttE8kMrBsSvN3RuetJzLlwaFLPn0GH7/ZG9ZlNacxHzmn1xyAkhbhW8hy2
Vj6U9dlUj04L/3gofm6o9OJHIaJP3MMEzmtw8fxUb1Gb6EJYMy+5Wn6LXfYZIlTYgrUDu9kfFP8q
Stdj66uCZdMMVYqJcCtNZbLdG0Gs9fDfMSHeziIndq8J+0rsYVP/k+b201m2X/xaq35m5ARNHxO4
u9Zs5jdvb7DCSnVg0+eQPph+etv03fiuQcVyctBN8j6lh51GAgwX7elmd+6HFRLixY6smn8Desi8
A0NWAabPiVyl8G6KjOJT0dOHFKOxFirNS0rB29P9/gPfRKGNWmPRFvScqYkFgejkmOXu7StO+uOO
cYybd+0EOO/4bDzbJQ3NOxI7+aPb1u8Y+RID+P04LBMeBsGUjhmkForXS/Z4CPlH1C5O6PAD3Smd
s5SvYxAKedb6OYM6Vcr4/dhxwEpLWF0c8xxILaYzfIsRwPNE+IuoWq17fDdZdZqjMqVbr+wXw/eF
bpLOceimRnlUP6Cb5LTul3BZFX2oY4hZBpJXhkVEVut+Rlf5jrewfP/JoUmR2Y9al+SRwOjOTXAs
JVlvXF7jvGxPqs1JtDYUiIrwc/muwYWFAOlUxsPwhGoTbyFPm+2TZuPRfCP3u/r7Cbl5nJzfaP3f
WNzfGaRr3G/Mx4SpZmHe5K0dlKQmxB8H8ba9r29ye4M2+huOSwWHIougS5p7DZeB8DSmnpEK9O2T
e9ThOaaOiXusZojCv79+pR02Km47zQHT5y6ygQoJhSyWLEFFxlfXI33aMejB4Cmm3bbr3nt/ApjG
ZF4zXbatYQHY+jM7YmdW8T9JLxWYFuLN4VFsL+TIzsz5BnPn1uCpz5f2yXUgJnhHs2y1+5F8uq5N
+Sh42dazHbaBXh7/jxQxQaI50zajJbr1aua0+EB6f8wogzv/+DsSq0GPSN+GN8sxwyK1tCgGNuMt
Y+QW2dADlZ4eVNw1+mG4ZJR2WtQsxD/MitlI+VoTaBk+cSx8z/47aFquvvj7FEk+t4ymqkKxbMeF
xoEIkN65+8RXpliNnBaIr5sRvO+FN+lVButZWiQBbY13QBq7KiQq/FYAvORRCuH9kT6+jY4Q5Ip2
GLDPbwfBLKNc/7/HslE7bI9IW57VYSIXp2dWs8V9kcm7bm0ex5oRLcoQNp9fa+hdMYWrDVeFkNa0
i6hDdGZUVSQQBataZtL1oZH4UUi3tW7p5I7LfYMHFB7MuVUB0A5gVb3jJNyhqyFjH95fZJqnTuDP
oWtKyV/aGccrvq1yw88yWBb0DqyHgn52OI8bh02iCQbYLDlF3Td1A2Fd8JP0jPGRwx5UrjDW9VC8
+9SMZyy/aCrDInbXRO1QDQZ1qCdhWloemny6GBm9KPBP8ekbJtvZ2CiD/TQQH4UnFIinysAdp45d
j4YxHvBieVL6NRG2xBpRAxTRSuhS0bFY+jgpi56yZRBQAkHrj7WVIkpAen0KuGq1BBMRKHYT9VQ4
zMEGbiO588bNd8bY0N4E9LNM8/rRDMPkcAHmTLUURZQDDCJeFD6uFcwCh5TYu0bZ6lP/UKwDll+Z
SdmuZVDJnXlx3Mww7g14/i5A8Qd4FJXyofcAZu4dhULs1p4LfjB9uWoTYplj7VthbjsClD+3beSS
PVEFNIEqbsSOupnQTgrMY3vjgPEjBUCg4zEegtCaafUCLvDx3j2UJSBMOYk8E490Apcr7V7I5nFF
QhWAiLChdYvml98thzHbAJhhycCXIZdjayNVCEzlNY9qSjB4FcfVi7yCCq0cJB20f15L7Wf3JZG7
kCIvst9XI6vaNHJfpMf6KyhT2SG4M4PNMLlWsDT2C5t2QRMzWEhtJm2nol+qSxZ15+O5n3+pyhV+
oKKj+k04YZokTt5pXM4SQfPqDnxqPi9KcLoDso/EJjjFsGOPTfsjo5BVazwE0JYfv6eKs2a9WTNl
HgT1cHf5gFLzzUI6h6HbCTUq42CU0s5yKoNyMfPlfN2uRdZv8Q22eViGKm2oRzUpc7VFaRCTgF80
+/XG9tkaPhaY1xYlZSTuvnVNegMXmXD8LiPwhRjO+9m0edUU1Oi7MG8/4yP2sVuvFSqJf60qCHcq
dosA1DANO4x2u7QizimaeN/+b9zjXgk6Qa7bdMonzKmIqjMdEei7kcJoIr6f9uwYI5Q2LTlqe7f6
gQeGiP4MrlJem5RBKU8PU/TjjY0tYcU8ghI4JFR7PnjFbl3Q65qIQ775Ot5z3Ec8CjmB3ahtIFEE
gMtnS0ZCoSxLSZOK4JSShW8zOg63GtBdwR/NFq7OUgCNsFrdi2d/1xW9JfC8ABZY8QTRDfx3LqWM
MWA6tiOBHLrzeVxImNhyrNTnz9U8BbEg52w75VnoaPG/VEuYaIXjzGhynBVT21T1eVgJ+Pz5kv/S
w6DlRwbWLXxfS1afpfX4+bGjtze/tsU48TJEJUYL6snHE3Bd3JImPIvW6tOTKPvgVnLyNwDG4TGP
QIeslfiE1/T7Ya5g66jZz/KNRlB2P0w1H52XYLLt+kRn/kHU2SrTjcPlyXJsl4l8K09MkKQr/dt1
Id/tQS5ymoIVi+/FJHCQuYeyFzEMNRsAkj/JAJHg96CnQyWZc+ypucHC+NEeGbL6prT2fwzKTVmS
PasjeXyQ+NJnnG6a82hztjOfINdNynRuplBms6+3nGmoqz+/+EDwWrMJx+CxaSUYSzDjVOl574dx
KLYDXtu4YgPjik2jF8YLxaEp8iXbWAA8/2E9wgDxtOKfklty/JEERpE17XlrvzJdrONUzt5DHzao
1z+it0fAGtxFXZRcc87vL40j7SdAcm4OCKnnXSJcrIoOGbvpB0KT8RWkMXODDDfgunoDojBgyhD8
ZiiFLCR7R1Nlvdv4QQzsOsTSqd0VD1z14GMLtakLMipAw0d97t1R/PsDEMn9/9Tjy/YHwylDYGIu
S0sdIjlaV84cgowOwsm2t+MZRYGp5Ahhs+texaImGb8IRdtr0bKBIL0MAv7hqRLli/RKhO/S297W
pXeRp9xIAkq34BieTq5I/OSqrYjtoY9malnijr916Y0/6NCxURYhXU66RWBdZHqwkICN1f9zgbHt
qK4ldVx34W67wH7tB09WA+zkivoGm+5qwIMP7nthBJ6pV0aFDkDIt0SbsRzNyG5qvCHse2gcyRUm
R+j9CaSX5MmQx0QTFX2y697+YpvWSzbId4/ihpy1PmB+Djj3aXDsOHMEGt3bxFWYXhRSXKIN4oM7
KrOrmcQ6i1t9fKFkNTMuAKGEbz03gFc0GBFK1VikWRsLRPfuoUY60RSuwtM6KBQb+Sevj1uy2bMk
1QY/cQCjKtnJWYVL3NAcvgy6EohmJ1jR3+AO/DhmfMz5OgruCX1LLmEsaiTM7Mjjbgul52uSzBuj
xJZawSg7TQ4qD+5nDb8f49+ZFPGezhGLjOY4HHiH4P5e3QJg32H7+c6QHFv57lLZHoDeyvFrzbcc
tSI/cckxZUKndDaOk92woWn3eQIZjcMakRvA9d7FZzm1eXSaDISXhplYCyrK3lHomGpAyjql5AVv
CPZS/kwvP2kWxZzkQw9e3esfxWT2tHX1NsmLb6VajIqOYzu8uJC/KRhkTj96hhgssoi18+4vcDni
oC2uv9NP3Jy233dgBLifra8qz7F0daM8iRyVHZ88uEoabhHSyh5zdVM1UGyKzlIJHhRMNVkttXeq
mpZdJ87cFqFOhMfAYj5BPFLl1A+lAqT2sr4pybqE9U24tWn2C3XO6XkM7Y0wlPIMsg5FS61L4AX4
IhN7o4C3Qeb9l9Zbt5c4Tbx9woHt7LGCbrhjNplAgUNHFrpdd0nkUUufWRiqnr/b4Gz0KTrIm5ga
W4NHIRgV4XRXByvMWYHobayWaq53aWhTYno+AQRZZs3BdTUSvSmDdvE41OUp8DLObNbk85jI677G
o13tBdcdcijlzGAlM01GNWQMgOpH7LBrjt/Zq5OBjmviFCy1YN+RIjZYfGbcJ4gpySBBizI44Q9u
dR4N7BefVpbLAGPO2H5CQcrm6n61TpIH0jvrXbWuMpafaqVDQI7YLQ8zKvGXnH6fornKRgQJehAq
AlNKMf72TWtS7Q881vxkFFAhpDYd5FJB7cnL1Fo14ABT/uMlHkNebBCFSh/S36Av6wx6ZsDXXJnq
Nyw3+NSPWqVJZeAo0Nf7Vv0jj1Fzy9+lcQZVCEAWokBEkbLLVl5GWCpvywPDbDYlNbqonlAHx4Lq
OTStVyr4gw2RPoxQrth/M6KjC9UoprshvvbGx0ksrvy7kJgl/C04teE7i04IwMb3ndnhTbSdQj4d
aUUnfisLU+g8x8aOaVDhCnoSZ3stogF228UfDGH3s7jDKhqiS/jtrbyYPa4g1d4lyX7xzU1e8b0z
0dpT0NaG5h7xbPTdoUjIJwhQ5O2RXJtCnJvIT9szmP5HUCXUTlKesPF6obk7UI4zfS8+bgj8EYFM
omAqhaBp6R4nbrCdsLo3YNkv6sAVYaulTWpTExZWv4KCpqrutwvRwK2RGEFT0WqhMBjEabBmeYCf
Scv7x+P4jT9izwVMHpB2FDUrg9F0fYKKMikNDFWTwRHRbM3Ky1us5dHLGWmGW9+GvoZfh5z9wK/D
baFpiUWc7EOtKELfYswGeIcXvStbt94IGhXpoU07J2jPORIS1WrLim14kxlLaYmWHHJzxxy1Kex5
9NxJj/CVdA0+EcFh8DqGcCmzKP2WieG/6Cv5d27+PR0cmDUs3pMTlmLbriw4z4S8RsxxYop0ha7y
XU1DfA1BOfp5xetXg+q4pVX1Se1GAn59GJU7WrBXM+cJhej/tCz0dKXf5M1JWzP7JH6QxJRZ2U+8
2VqxrZFtMuvlXqk7fXOGSEAUAuPIBbHIWGyEIycn+wyXOY7xLjTDFpr15lGFVUe1VoUtPaOAAC6y
11ByMPs8Jq1DvpbCFrqcb91n5FlGIRjzsBozy0ZMuc0yr8dVqIk+Zx38ZygqeeTOcUielDI5Sf/9
NnE7S5WvFDlmhIZrxFQsHgeyV+p1GgkpwVjJdRKqUja/Tw/fny+F5xTPEOuzE9pxRqweYBPV4SHg
m63mq0r5xgKwEr4VvzCfuQrkqk8xgewrCHJredAvZniVaFgsg+BhY6/EdRiamxTGtOZ6UFr6dw0p
pkpzlSCzUMoWHPNfHafucTHc1AqEMYsR7BdCO1YLcatFcwl0sDm1VZvuhsb6QM74EIPEAHIfpXQ4
18F7Y1ShS76dka3Jc744ZK++DR9SFbq6vFvJdBMQkbOzhiyibr0H43Ho2NDLuqESMDoHAV7tEw0G
zyUXFX2syOm+rDWbkyqBv5wR8l2uyaXq3lsJDzGOOASmDPFjrUF49BzyQU8U34OzOqA8rp7Hppsm
qksgcwSURzmr8LF7ujmUeauWlskv1NF2y2kUG1hFEppcpzP6wvlycWitDAHPrjGtcBOlWfspOD0k
75Zj3CG6LcI00K8wGrKW4eaPGTW00A7m/HPEboet5kCLK538y0ZAzS9JRwIYPXbnZQWFdR9Cz2U+
Y2sdmTf+IQK1sSbXwKOu+GoGNUNTul3Z6IHWJXNIWfOrRzeKrwZ56zlYISTrBIbFH8MXvlanjk9r
tTO+l3j5crt3kyHh6nXuntYe1v7xwdx4dt2V4nb+/amLDM8Rkuy6Tp6TNEGP3M4ZhMwLU4EvscX2
5IhUUzXCrpQTOdcEXG7RVGZp2pgMpzWzvJl2XU7Q3l7P3sZlQEw9j/Pi3TPW84qhRT8so552xlpd
KsFjhOwxQTFfqybgHHuUPR6nzNv8OxixGtusA1nMgkbs6+6LaPUab21XblLChhJQ+hPwHd0Lhmcw
u/wkTNMOMinAAlewOEzZ6uFkFUzWRKhng73F9VvwfjKVNzT1aeWLrPSbopn0PCtIONTFAdUDuX3p
i8Jb2Fu6PGmtXNUMbloF39N2TXDU5vVdsaQdSMFU7dV8+pXO1pKh5mElo8suQ5atBb6VfU+xwQ2H
rz5g4jrGfmyu4jLSP0Fp6VWLDqS7z4vf4kz9BY4bI7jDj3Z/fxufEaSczll5YqwJHV6H3+JbF3+D
gvIhWwZsvp62ToDPGKcNhYCCfb7+Hnj3jNz+lvP6VJdAkQSuBlfawv5fZy81SX7ohgjyBerhZz9K
0uudyGfIujw8TcyCdt3ixsl/hyiHfAhsJYyIYeloFNvcpzW/kCEHxmBlU8yEcfE8+5x53aJs8AG5
oXrxuhIVkdfNd1jTTYbZ/savuTZ0vqkrmyrrn9jbdkQc7FdJlODjcNc4Q28ezlYV+Fm8ONRM8kil
3SGS0o3gN/KRIzAjW4t0dl74RF4XF53TZ1M6EldtLWTHZMytlNvDj+fpaSSlz82P5Jo87vqGtNTj
7E5N4fyagLtflQ6eZHgDzu3E3Ee56TCxD47bz5FsvayHZ5YELk9BJw7xevm1ZWSJckjQkXg0F9C/
GrMoSKj/pH+c0sNFBXFhRX07l431M0JLsRQnD6fKQedQW8iRbgg5D5voyP0Lehc0koF0xZdcLV1p
Pi7Mo3E/DCo3tvJ9O7pK25srhO2CGi43duqvxUAMMX2eJ2In97PbqNEAksI+OjvizOR9Ov0XjjPw
UFlAo5K6a/k83ZDe4ZnZ9NIa2Nq3E42XRbhVDJm5T6nujd3IKDrwyQQ9njkk50LdD8EAAlY/DIoh
YJhJ+wGMNufNvAsmCxqA+X8Jr1WcesYB0LIy+PTG3J/HN2Buxs9TWOxZkwveJ4ZowLIG0/jbsD6l
dFFbEynfjUhrHnqBsqB0zpoDzXXBj8XkRVfhHYzqUgx3LzkcQmzK6JA83Mgd0OYJXHklY7A4V5Gl
gOp6+zAxp1zFPiWY/eu2E2WPQAmgDXcP2D38m7s2q8gxgjlR14ZvkH3Y05XjvgnrrHQSYii6NYHx
F8rd23fBSqU3AgrZ3S1tGB6O8DxhurckQlLCZK2NNQkaDT2xlCaItDibHF/VZCL6dsU7xdURgpNb
TXMdNpmyG9pwUTPJQs9TKsd0Ot+yh72ThCvmB6A0jutyMBDRivS5MT8arHPfzpIGeQ3bmo+pjU/W
0fUBGefiz4upEYqSJ7u1XElXv/IvRxbpkUN4nU2PPVQTDsTfKT+ovSaBpd++hihUX/1zpJkDxarT
uib4zYZHS59VWSalm58vFYEiWExvjT6g+vuZSCS4ZBJuZEO1dBerAD9qeELhf4u3linqOlXc3U2a
eH6lnaXXzcWFvZJ9ifh+jeN4Z8R1CJWmY5BEdJJFRnQ=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity ps2_fifo is
port(
  Data :  in std_logic_vector(6 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(6 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end ps2_fifo;
architecture beh of ps2_fifo is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~fifo_sc_hs.ps2_fifo\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(6 downto 0);
  Full: out std_logic;
  Empty: out std_logic;
  Q : out std_logic_vector(6 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.ps2_fifo\
port map(
  Clk => Clk,
  Reset => Reset,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(6 downto 0) => Data(6 downto 0),
  Full => Full,
  Empty => Empty,
  Q(6 downto 0) => Q(6 downto 0));
end beh;
