--
--Written by GowinSynthesis
--Tool Version "V1.9.9.02"
--Fri May 31 15:50:54 2024

--Source file index table:
--file0 "\C:/working/_Tang_nano/_cores/ps2_fifo/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\C:/working/_Tang_nano/_cores/ps2_fifo/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.9.02_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\C:/Gowin/Gowin_V1.9.9.02_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
t5uPMPBn9HdXo3+vH+z4h8vOPjgnIL5ts4ZCADIUIUq/luB1tC29RTYVwtWt9DK5RvyPNO/1U06/
Y8oJCw/CqVqNmQRBOac8UV5N/rUI40mxLIRIvk6JdLJ15mstLWM6jQsm5p4gB9qSxIGarLMwa6Ze
HZVWJDJkTQrzA/nz3fpDnbG6QlOPLbASNSiNBFoTVoiNqe4sIa/DllFUPvqYCTh6cNfGzslQxZmu
SJ7TbhUV4RbMsMNuH6erjhgWLpxSXzrR++uj+Wpj2SZU/+nqCUmSeFQwNovegKn6ogSACnf6bJK3
eoNiWn4UWPK8bAffpXVNACpEwqu0o747Z0wD3Q==

`protect encoding=(enctype="base64", line_length=76, bytes=11168)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
FDXTKAtxAjNjO2f6bzJ4JzmM9HFWv+B4qS9/R6ubOyd8ouKmGNK7JHCnkHxJZoz6Rzztw+Tvp0Og
VYelhMJ9W+GsKUIxIP3/wV4SfZqkK17vM04cOxa3CFYZMrvocEr+38rzsvy4lyinvpluZ60XtctH
D6Qqg7qxEOI4dWpquA27quosVKnwYHecvNRbvaqNYC2Cht+BE2sa8VeBb1Y3CjqJYSWUKXb7JSAm
WpSgfefNEB6XOa9oZhpmn0DVyiqCk7eKn3veHtDGPZ/eak8nwl3jy/zSpSAi1IZYcqwOgxEgnsPr
pfvcTbE7ESFL7y0HM6I8I8BaAt8PibycRGDUfsWMJjHtnX7zhp04RV01rcq85+OkOky+Os+fM9uJ
WMXJr1MOKQeOAtmKcDDrhA8CwB3mGkv7OjRxrQgkXeEd7Rz0FEgxW8m00rJWdd87X9VpP6/Swr9a
ZvQxB/aM9MgkDL9pJLwwSWfP5nX7i/giBBkd4q1FwztNQzEIGXXem2rdNRFReePsFf0BVwviyXt/
DogRTiISqH4pVhvDpBRHDzbGuSwpWBldnqRZeqNGOYXmyccovpLsRSppiRuis5kj72lFPPdG6lPv
gHYlnYTvTZIm1OaK13qmGvc+EzZ52MlSFHa2PvYaXWivY/Y6E1LdontRDBbWEwqutl2yRS3TqIQq
sH2Q9BD9nlcbVE6AB/d3EsAOh68QwnCpKS9+5CLKaQWXoS1aKifTCQreImcgyqCHR4/h4iS4EET5
xzdnalMdpWXV5QJZn5kECshmIPVB7gZHrGIRW3e03KlVjtvvw1Vm5THyUjyAnRXkdOa4jAZ9diZh
yl9DekoEx2J2W964oDBpEkZ6F5nDthuDc3l7fSzvCvS+LRmQRWJeAy445CQIaGo5csIycKCh2+Tk
Ma87Be1zVGehlfWVvvwUpmgVJTOd8GUWrx957IsKrjWxHaFxchJZsyO6nC6k76c/LcBKWlPUEZqL
x6j1hAxLx1ePFlqOzAkk85lX6iU6D1BfRjYCCQUBy/Ab+GUubWn9rfBkd4YyQ8FeoS+6vWq1MzeX
2arN25C921ytV/dA/ymXbEO12erxmYdCmTAJIe1dJdFcAtZ1icvQM4RGX7rWFJHU1ug44Nl7oCEm
AEgJ9+xPIxnQZ955Cv/lhx4bh9l9OmNdUC2uHlGycrV1+VzbriFkKvCBuplhMx1FZhomlHIWiN/U
TvEzHnOQZc1aLJRFZfG4yEfDYhXZ9A3y2giZn8NRoJoYHMBG+pjNH3ijQ+SVUmsiu7q5iseHUCL/
Hina/V10UcdbJXIOKlEarIT/H6gYSAT2aVYyH9jemRFk7PPrXtTM4fozFzsgjaAtQLKtOkUbGCi7
aq47wmGT5N9hPZy0lYpH5iPT/Ekn5ouX160qIYB2jQm/Aq3SgU4tjF4Il9L4J1M5v6UYVdXPgkyQ
urmTut4X8snhCpiXzvzVYchVOZskqH7YDWJN9MjkPKk3IkjjKPehq4t8lC8PpDeGjwgcbmN1G21u
9vtvFCA3hfQxef6yLx69zAXLg5MB7O/UthcJoEZDLtEEKGlo37K2D6g9csOY3KmB7tIVeQsrZ1Hz
lhoXGE5Zf8ikVT3ybegWaxf1eb9/LO3JSiXF8Mc2CLRPULBT0Kd4NTsztKSeNWaQG3tIU6rV0xol
O/X8I8ufAH4285TDtYcwNxRLy3je0C2JJsvsBKNMrDDBE27oxChqomISqDPf7LkTckGtDwKn1XZi
mCQCHnzPuqm4bxxXniWFXqJUkKtSGD/1aKsshq8w9FG7gr/OePmJPZwNnJneKh8+pPYtAc9Jgafp
+psO1z++BeoFrkCXlJ9pam4aWlB14HbWS8TcdbqM2AP/tZE7bUUafYcPXa8oshMeLfQ4GTc6IYIi
nb79yD6HVi0Ak8bM9pR8ECoRNoDla4QRqLcqaIMSQmkd9cN0Ka+3qUMhAuVHfSXqhEtRZKmKtmG4
oNxLZeZPdW7jltijVIS7SyOd0nZ8Ro2lLHZSWs0srcJ5HYi7hJdXHQw17u3VM/XRTDwWXC2QFAjQ
G+3GW1b4BDYbUFBmHcZATX6kefI2bAGioqHRpGw92TL0dX84kub2rcjC+uE92N6/C6I+UFatwUX7
r0nKIKLIUHtmzAfUkJQq/nKJxAxJo8sVlEltbh2CTG3Rubh1U8oOdnm22iHo1OOCemlsMM7tVl+J
eqvDe000mEIOptTniQoHQcVnAT6tVQ5FwMGUenrBccBd4l+3AW1sBHzTOY9JGmHocyex+0WnIQbR
V7a9Rjq9+nZOYBqmkkrQSWK2oIKJcr3CxGoIhTxgiXNy8P73SgpmLhO3VROVZYXg3xZCYRC3OBBG
JyTpgXLUzQMF31UdSclB0wEA8VsBBRgtc0bkxEU9LNlPbQ03Zvcn4g444UC49x+/s4e4mCr3Mgde
JuZHnCcwE/KXLa+TeFOa+dYs+tytyplgQ7kYypNZA2MshrfUXsB8OZ2s5WyfnCXTQkwrvDTnhET6
cQMOCp39CUrPRD5mRxwunoNSTWQ6N9YpjawrF9tEL1SjFQbg+TUiP+OqTqDdzXnVIGo9o+sk0eKo
uY3rKl/yjArCuGzCkK5PZwXoua2ADfN8wWHDWRfJj+E9+bu88utC6m4KvLAesfVeJUmfwdpzkERZ
Hhl5rELxdxNex564RzsVmrxGfX6wj+P5dNvaofjr+722POL06psYsTRDQmKYYF4RF5yxqUShD+eM
aSwj1QWkwRMj3DPoml0he6M+wqfXAIs0ojyO8rcFrrbBvRNWYptPH+mBYoCRDunvf1UviuzmFCV6
4Ldys7FLlS6Mxc6OtiBvLanlTz+GVCt7YE3wJrlx/G0Lk2m1zmFjhByAFat1PoLec2iQY+Ak39F/
9olRYgL2K1Pws/HZxY3Wht6YPQLlSOBkbWRXwo79YnqUMEYMJM3I/D06zTXBlSUlr4rZ/o/UY3WL
Wr6Io73js9gHlVb9vlBZcQB0LA2f3o+uUX/WTiGXnJ6IsrTtf2PiCNTmMp12wi/9FH8WvTXuBBST
4EvR5ciyQ5uVT4BOUr/Jz+p7kOa+An6fFXebT9HaJm8v38I1q8eeHZ+ck4h3632ukFkWHtQdok+R
SkapmWVnkzJa6xno/OeIWYVr2g1JOYJfbJM4Wt8WqgGr8/h89Wx7qwjK27FjE7gcF47IDwQChbHj
3ZaZbrdou8xf59h2ag7nwM6yh/7GMwkPTn/xWtrYyhnvw8YWmJCLiVShnJzZJNgazIxUKuJ5qFV3
dKVbSPstWTqx9nWZ/eLfDCoch5aeXbi2A5AduyImj19WweWg1Phpe3o/SB46r0qNEnGnU1SyWPoi
cAM3B0o42/wLsKiPk43aBMabn/T88oJes9Rue/kloui62vDByR8+7AiyXGd1Cd2Xr54KKhuPMlVZ
i2IwpR4ww7diLClQ29HEGt+CyBK2g3+m5HH8RSesRwixihwE5Ty6W9jQOmnPVWarWc7O2OH3h+Si
kXaI+XCbPkUol4HomF947V5Lz2kwp9YW77y2hSk9PoCfuBnh3PQhAxuwdBEbMgQefnPP68qc13OY
vvVAoVgOTS5BJkCwuiE6Ut3EfsNMbepOsgVDvtsKEvU3lVDFKSpil6sIPdA7azOwfNdoRmIt8Nym
6Sk7KE//M9jm/yYqQXS1v47Ew1GLoYSghaxJtOBNC3Yia0zrwOhgMEEasBxe3K/uJsdl63rslfIf
G3c/lUrCr/szwJnPcZjbu5ipd4/woOwbGxOdWX/7bIxfZVpo81mPEb3bTzbbgNX2WfNTV3riaFCq
CMh74KJf7pjUXilXB7XWTrB2210SFXAyBBTTM7tIYdN4hc/Twq90v4al8dM6gDsKyFuPquzb5/Kw
voMP4sbOjj0ehWkCXFIkdAtGcttQTx7n4dqLi6rHplzd3ZnKwLgFTjbrfJmLamJCi6yLScpkKLBQ
kG3piprv2vL64sP7BUl1K/ellXAdsyiBqE+iDHtxsjzYCoj+EvdfKjH8KqkXj0p1yy/wDOgeoKJt
OeSgH1ev2yRCuW8XH9MAggmKKFoGdofOEhoPHGDbo1AC2B/hMQdE09ASJmcYpFIwztPTk4HGnA9H
ft3o7E4jRwDU7C80qqZNBhQK8lgCQKizUSToFpgZ+bLfE2iM1QNotdpTzI0zK8nvS7fJy/X5oaWn
o98EIGsRg36lThEhnMaxdb4Y6pz7TFEOooQjiRtWYT4GAn9b0o6ZhguCy1u8w+026B6WOlmwiDc4
joDbEg149/oRHMGcotJ102+Hfu5r7GJkomVK3djUH5oNLHzgCM1/61vDFvlYBy4CBhoNkRgpLFEv
AMJDsLkKD70Ssq5TV40XzegbVtZBk5V9/xiN2q6+3CUNVr87VrZnNiynbi16gCzWX8okLM5KItE9
B7qTeEElji1SucDv201/j+foRPoLNBkR0B+mmZuptduTRG3Zi0Kf7oARcJz3nDXlaLj+umwACZiV
DgDbQR5YgaYY7VQgOm6pw+nKXFNMjY+bvZwjWI6yMcZE7/fqGkJKtUnwhySJh8087ZbRcVLcqhuq
cfny+GHzhWtWZrjDjZJA4OePg5lmWPU/+j98c2rnIQhaUjhOb6KGRuH6dGstlHUi12Pa+7QVfXlZ
WsY9lEoMcrIywxPxdwLQFKkHpKVPqd3Dafh0zuaa4fdN6vfIS1EC1yJgExr2gJwJwS1wrETfoZGc
gAcKP2x090P8TbT2uD31wDHO3W9ijJcLachJWwUkso/oTgqgluEc1Kd4oAmv67CxDJQWzi4BUtcn
+M12NjoSTWqOxn84nLdldgiPDYIuJ5CI8s0bXSNxPUBxS1ZEZyw0j7femGcfp4o95RbsPd+mF5yA
tmSVWyVGu/y6DoZErmz0GOekrPoZaSTIhkp48lxGjZY8tZ4OuoWvJiscKx6HoZwxv9zgZBiI/6Dr
Ot6sMH2YcLA5aZN8SvPpJJdeHBOJWDXwEDFd5FW/oPFsG3wtE/Ftb/o5RLqKqc1FS7mMIZrDryUN
gcHgS7syA+5KD0w8ugOk7zek06DxNAFEeBSEkX4BnFPmJ2SJLZrDkRvaGhnmMk6+Xytsb6j7A1+2
PYuGdQ/+LW51B+O9itqVsZrw4IKRSJwudahlPHNhR1ftGTKs1Kgu9yJRjdNY34VPfVsOplUBnRxU
BEcNZnUGsrk63fMGlzYE2uvcZGoGrNsONfgrtXntn7l780Z2ztomE5/6IMg/sy913l6guCd3E6jm
kaGV1cUIXlHJFnlzylt8G897KXXJjH9/xwTZdRWsQ2B4DSm3A6iuYGoq2bmYPEnGppECEc/2W5JK
SqHDfAOuZ3jkyPhvEBcPRX/jwz87MTuShNttFnMhlbhqFdL3ONDUFSKfiYM5XHRO/FNu8ArGsGbj
x8K6nde89qQsOKwrbPW0cqSRcyblRYGs94Crtq15whl292QAXuUegtHHqqxNFV4Uf5Px4gRO66IR
p5mnQAxshP5LDXOAHq2ia27+mMRGSlF++n8krRhMHTPRQeXGdJNH6obLGDhZlfqjfM1r7cSDTIzB
qyEQe6TdyQX0Ao/8MLsCoDpa4ALm53OOMIPdFzBUpd/LefcYGfQWwo8zUge6tSeZqfPvjO0PawW0
JNARphIXF9Es7jnnBSoafT/hzuBsG8XwG0jaaeZ84c6JvPsmICgZRh6m4tsaKf1wE6gWnT2r+01H
cGbSGiZbTZtoqYlawI4d6ICFSm1/x4WkDEytPOV0hMrBs+mbJPGX1uq1DnSCjWKl2djFUC/kOdPi
0XdJkcgCmVw61Y34THcUDuS7vljD5ax+IucgJxZcRXUDwqp8g40nz6gkvEWEF1RlVvAsjBs3ouB4
jYPLqF1ES5niVVb1TXYEW6RvSE6WnwEzCGLIy2GQhbztdhJojivGCzvgmwpeut3KuUIEtg+PVkMz
hFydUV/O4Ma2X8xt/Kdve693Ov+nGkk/gX2UhmAEcm+THPcJErRbdUKQMXjbkHY5Ig5nkuacqfdT
GStsatGxPnarzqEd5ExJG2kEy/Rbh1cdFwPcwC3CKkfcDiOWYEbCUMX+tRU+SNEQT/99LxB5TEnz
BA7iVEOwF3IynvBGunYBwCxvSo549AhVOqVeIEVHxZQW3Q0I1r5IL6au8hGLtgn90ndImdPhl5ID
t8G8upzxvgq679C9726HUJYGKRVoEC+RmYkZ9BmZVnuxlgm9eTSIJyTLIfikZYNQ54CSmc4mv1lq
Heb513AQt7SZumFo74yzVRhaePQnmNlL9oGV3K995+zYGWT1IkqJKSn2GjNTESbMi/yJN+zVvU8S
XSFlL+kWbLp7T4o6DPUVG4KcAlz1IXhaVjF8ZManLtMT8cNlYefWxtZ7zDGpV93n3RLTr+BM+gx7
pjyHJSA1cI4kVryx+ZrzG0l/rREgPOauBFcw90fG9mIe86rQRgSuM+COsAhr/FrXH3HRQiZyj3VH
kWq3AMIMeLCl6oSgbRdqrPZ+MNf7gCrhH/HBHd07j5P5rb8VDpjPeJn5ewjBKYFjsDWsl8Awm4vf
/WbQ7mNWeXHsbjYX33jP2dPYk325VJ9EA+vx4vb+ScoYL1GejKBxUMHpSIv+nKTjDS+AFjW66EGJ
ReQ5j026OHfr6CJSjajCYuQgKfz65KJRHKhkpgSvVr3EjGV9G0LyhVVC4ZAS99aDbVLurAWmhnTj
h2m30xelVklTyOKUXbENIY+3HJmqun87/rt0uTLfaEQj1BOEXCqREEnwMwblOMonM0Cm3FhMVcmn
wIP7WDPE4NySNGjjxAg3Lp9U9aGP++m7oDp4XHmC33Sc7AdkGDJKl4XORa6t0jlBYgUsNUqbixpA
elGui50Jn+7eQr5f+IptkInhJ09zW87vFjANrTbGTQ86XmzvhA22YF5e5h5kmigIG1rppVQsvEZ8
dWLs4ywMVWdrQBybMLlPlcvvDRqozL2ZNuJGr5VONT0tvVcJ76pIgta4qj6OciGhE+4BrUcEfRMD
vLbqfbzSkDk6Pst38865ngDSCaD9OGJi2CbirjtkLxs+LmySix3YAV1b1nBrn0BDW9JqExxtsLwW
3ho69rKNDnJYT1gel1E7UJOcMb1huo8u4aSPkAJy2zzE/rKcB8MhXaJudP5XMU1mjMGklSfZHllI
fTGuvvQQPqD/GXVBpghn65ISqvdC5z4DX7gQKrDScao3Y7GpOlXfSHsruRMZFUFqelLuQLZjYQS4
3fWdo4rscSRiyjJczyc4hy64AVE33Exb2PwdMx3pGbQaoIRcJrsqtIZXQkJXMydVEJYgYa93ZxF2
/sY9SbwWFBDJ3kaW8+5OhpXx+6evtPGJKggb8gAeP8zFWlOQKpV79fT2JCIT7bDQidsT4HfLx7sm
d9eqnoSraJtIFdRybXZsd6fyzo28FWlINsxUSkBn4QsG7E7B9Q/7ZuP10mqJrA+3fxqrVId9X6AS
VQNNeoXm9HWqMX5mRQdrw0PWmHMVHbGCRfgP1k2o5afsPdguAMbn4uJsw83QeVvRzxvLetbxrgYm
dnQ4ePIEliMU3nVhW+8rfeza4eQVt40z7cPfoiVHcPzWskZGY+s5+HRFvjYIuVn9Nj0aByp/K/UG
cZFBS/qyMCUCtdtxT2GrJ/bXqNsMAIgdH16vFxJEZApOsBYK8pex15kBmeMCTpu4QHuCnAhof93B
KYADoxm2hJ7zqEs+9SoEkQO2YIQQxJtFy0AiKnrWXCg75RqEVfIQeHONkpieYrDOp2RnK6IMvfik
PqC5SY9sKLO2yAUECraPSEVd+TeX8puPe2NR8+PAc63jGAze0+oHRJsxwpQg2VO0SwyF9s6Cuujf
AsI3MkirnSnOU7oBRQDunfHb2tHa+XF4NzDwuCxN/410wam1dtqoY35UsHDI5TrpPsv2CQJznfZU
LvLnUZpyCL+POy9fihgU7eirEytabww2pEMssRz/kskKH5O/iGIeer2pVztD9Z3H3aaW+wNJR85M
YAPC39af0A4DbRiArU+UOs52S354T9GG1yBIq8eMA1G8KvZYev4TjtlnntaU2OKNSpnpwW08sv+H
+iK0gq89qRHPR0YR4VJJNXqskbz7hWAFt0dJDxMh93Dux3Cb6ckmNbo0ACEecMtkq/UbwanFeP69
wvcZdvKctyQUJfTHTjujV8BY6rEmubdp7oNzsM0OOqEg1JrusudZH/nZAffe1FGPIEigEaCWme88
pmvGUBbhYwgXKzYVPRn53fk32BctWRqfXBkh5CuehEW/o+gScpsMTzsqIDoqFdHmhDTGcWcsbR4z
YXYSwRd+b+xwsWc1G7W1gjXjz0+EkkKEwjOHqF/m6jLlzuGNfVuUgTdahNU6UhBDGRY4tO/Q4bRf
wXxDTVM4N82D3o3SuAZ8HcBljM9eFkLt4pxiWhDDgwTOUpbxeQ2v2z0VO6SGFzL5liyNbuUZCbn5
GXeU4aT3VSlhxz2N/mDL90bdwQMZbGJf/hvOtbMcVgJfchDboRSkERzgspLiktL1KMm8XEwRERxm
kS7Y3yZbsLFxA1kS26yi5rqPHkZp2h4Clwj9miCttwIFH5IMBs8OrpdPEMCy9IHAgcdUcI3jYx/9
7XhPFgLuV2TjxUCqkgj49phK7gHDOIfRDoU9uF61y7TtmUiFM+LD+wPyFU46w2Irgdlwmam/My+d
nA12zwvdG9dXyMh1IZWWSIs2uQ7STvdxIbQ47BVWawenry75+GzQNdZsv1SMQK2Fy8r8FnukSYdA
9Sx1iu8WMNeifQcc9bMpb5f6KbZco+atmJOtt/+d20i2VeS14raq88wfttbL3BSMMQaEZTWTaPft
86Hi7C/6xQfmtkQUBB8gaqzJlrEmw1Tz2QOLcB7wtTBz3chmCqWfg7gw5buZqggPKyQtHVVehAuc
/tCxRK/VBMrxuqgys/CZ96hJ87G6zzFO1agmTnNFcVL2ayZ9HRcao+z3FcRKPBDGBd1Y/Ef08WQg
jtjTPDeeSjZOILTcKJWBssnMHL1fwObdQwiVfz2C0wabaMq4nRXbaVz+Aqecc2RZ6AOv//wOd+4J
zp+pEzccEG+RdOfLYxLWMR7KvYD+LCsOaEINLjl3FrMKQ9SZVlFA48qgU+geXetYVRgi5B05X6oL
zjrwofLCJimL5J1P2yHJmEJ8NkCjk7w0/FUeUpkCaZaCqqyzsOJhn+Su0lWfX2LSGb0Am5Uid+08
sLoANKjjgFl785hj6BTA69u5cyHwZn2hM913OtC+RELJFv9tZkKraVOh4KIct/pV61ukSda4+a9+
dkhgb8Rivqnw1FfmK2ADA8yGVYEoqcoRWV8xTsTFy7TL1VJU9BZ/A511PYFBMHjfndJJUjtLcRM/
kYdBNvoBSwdQ9/Uqxs4lz8zUXGONdrHEojeeMfHprvs4KTY5Hsb3b4c1r8rWl/TvrafmZxLBDOSm
JEM5SvCGi9nC3lbXP+E8AGtRwSbrsaMwIY7RNQGTTrMHOncHLx8L4kpb+RFg5U/1wZ7KfJnP+oN7
FcO3gaQ5os+CQUDMS3Z4jD4vy9AHEyR6jKyL6tElxoVhlPQwjJyCaL7pbHbjcpOVbn2/AMo9JYUI
WGnRHc/5JgKbE5bT2Pk1hp/QQU7dnOJyW4PhJ2UC6ZPo2jc/7xxBgudTifCbPyiyIqHxv1WJ08B0
GJe/xJS1swvOayEa0NhFAfCp8fqyJjgYpqCKLjwgwg9ykuMvt0inxDuVSaOImvJdqQs3pQgYhwKr
fAQQ6xV8rC5vEV9siC9/rjXYkyItdM9cC94r5Gyl4anj0AIqYc03IZIJD6NjzUwvh5EiOUGGZlFU
P2CfV3LVga5AphSEJdrMps9ae8q44MImuoh+AebX+WSRHQM5/ddVncjJz60RDFy8e72bk1T7LMSg
T/pUG63mQDJdczDsgBQr6u9rRrdvz4eeb35D1Gi5wnV1N5gkpJkeHAJOR0L8eny9f92LFIQgC0Cw
ofYXQXXw3/EFMCWoOPi+CFPQnTAysWhY26ak0QXiGxRCsMc122XgOs4cOGOO5svxWzeT/KZ2QeDe
YVtq/Y70To/GtjY8IOidGnVh6r2pBdoHZ49HFfU0gJH2OFdFAQ6we4iYwcFoXVdyaQimS539MKcl
dejKSN86A9fQEvTfYKN2YdXclkmLdQ1mnKOGDNoPoUS5ZYjtlKksF2ZQCV/ePtFav+v2iiIJdZWQ
YRs/f+vMwAejjoE4QRAZim3UQFL+G5SOalZ1b1XWt/zHwbqK9rXBYTTutHvHz5VcQWgzGgBM6hzq
MqPSvA2ImtYk56bAYhXsjZc9Bjr3Z6hvsolO8e0/OdDZQaUZcIjYLw9C/3cNIEU70E0LEHsp0Don
1SPDG4PhYogmuNAFS4hkxmo6jMuSItzWHyTy1WgyPB/yS+5cYG8vYSiGdGzU4tL/NEQhlig9IsTi
24mIgq7iI3zyQvJso3o2zoNMek6aYMFvPmCXdalcumnSESAAblq66ldwSKlfFyJdRG2cMrDmNS+2
WrIVlcBmCbJrnbeoWw7j2xuNCkbwUnbNl7/Mqw2p9ARnwveMjX9wI+xNuv68jXXa/pSNFkZzM6G5
w2vj4CPOzneabb7gtk+eJw+5R5UyPhY7C7QXoyvDuJOokgsDRh2v1l8EjXvvtp2xJy6Z5GH02b1i
CFDAmkw2ugsuGFHMrnO1To1pxeCi8gUFcqeRB2oWB4pYcSnY8GWtsBR1J5T8JFQiXah7TFqEsSt2
yY0CDlvMFhn/3OhLMW95I5QuzBBwJZyctb6r2z1jSn+d3YLIn2PzEN3o0xonm3P7nmm5pv2KFXP4
PwBWVIIYIer96M2eRC7iUvycd+AyMdqxqc4AS3wyHWYJYSX1/Z9uA5xZx+dlbKItRzGKg1cjnq8D
z5Ysgaenei2StE55xtK9S8L1BTT+kqH/97139E5cl0G90yUXrFMxycYTo4aP/H4xiLgUvtZdEEIZ
ZJqOalYJUfRYOQKSMu76EXL0+DldQb2E+NklfyF/Fc4/oHMYejh9fxJsxShFekPxIDzocPXB/Keg
dkhYUV9zniZVJgwR5qtda1KTTZ906mhXaj8AsH26b26sUnNebL2rOOXu34e0KlKC5yZT+1EO6GnQ
FRYgjFVSt3XOPR0lP7R6mVd+Qh2NASjqhltmhDm4uDkpeew2EJUSabmNIpHSxO2aUB12JQyim2hc
w6ZCy8MxTt9XVPSdpEWgOjJDLiPlUrTSEdBP5Hhq6eTTL9fvZpUCK37utKo2mXcNN32dcOrRg8Pe
R7zK5aeF9S8bjK8QBXiRQqsiB0ncHevY2kIDfpouEnsr5f2e6N1bTp5+LswmTGwisgzlqmtk0Z9Y
zM05vxhTM1uGpKiZYF6tX29ODSquHg1IF7dywR5TmX0w08/j8jj4c/oOq3HgvPw7+VWvXQiJlQIO
kLqCAEYJsUPWZSysnUsUIXP45iOAQe2Oq3Kxq4vP7bgkYlgafwEh2RSXg+d21IhDk3t03n1YG1tT
KG3nFi5GjfoaG0Oez8IajGABAnGz2Nj8RMZfVcnjBdvtH6QyqmnSydXX4LRLDi37/Qt6JiYed4gk
TuOspiuv0lpzeuzJjiVbvR3B12BNslH6ELTCofB9JZc24Vq0epk49D9fqp5PsIBz98YolwxrOsy1
IKQpXRklb4c1qQjS7z2cwu4PAtujN55D3MVIWHC7UEKDkL6OU6a1O1iqcU2KYoQzpcpeEId/QwPr
Md+iPtJlHbI7Ix7Hije4XH23n/qOYiAfS4ArTNno4UriReXB5j+lQZqrxDOuhmGPv1vITiFk1dGW
Jpu28OrRX6vs7mr+oMlTmFRJpbh1kodlDRhQvFhMyBSi/U31vef8gjEbTq8azWjZsvZmsC3bzYuN
RYTrqfyky2NxE8qfMinzwAc4XZ91o3Xvda2cOzT5kkNxmGFBPYOBGPubBltK6k4KN+VZmlpE2v6B
QidZujDpvSh16D49sk+so4V1ugB/iYRkmEhVQBhu0s9OQuICSoC2Z8mDLcA5zxO2g/aU1fMk3IQY
w83Nm7bOOJ/4Pr2hQX0rTFLbJFQifPYrAw1+vfuCOSff8YmXNgDcHu6hLp0dggvBMdrQOjQlzHBH
vkB8awKW3V7DTFL/+GmRkCVKLJJM8cv7Xb80Chv92r1GF0VMa/iIHAvNUi1KwsXdDbwngAGZSfWn
Vow4yxL5SRPqXRU07Pm/uf3jUsz0zyZlyy+n+RkAfoQdzFDSjE+/UgJIxhAMuwsyuJ8LSGTp4AUE
7WjCU2KFvWwwoHT5GTO4gbTWnvb4sFJE9dZEQaLj+MUA/mYBT3mDQcB5uIJVHXJXOYrLCjMhojhc
A/NOVP6y3StFOzenpbmDMqGuY6zer2kivfor0nbDr9FLxnLKFIOvGFwenRmYi+Fn5IMjLdGHnKlU
GMgEqlXKq2ihNvihhXRMzkvXmMR1Y2q68S6UOOsSpUCaQBPGcORSzKDl9Y4exzrSgyfQzs49EUjL
/hB7nx9AWD0FIuantYHZUbQf55Pi+okknwFhQxg78cP9bZbF2xPhI6GNF51RcxoeMR4mrtdSB/f7
lo8Kot5Ql7DEjAtfVp2irgEYLg/L5Z+yg4F4PWJ+zXOWuvX/yfh3rOgPjIxkAqHFTrvWnSqNBDsg
ts4WYjd98IDWIm2DuP342deKL6dsF+rPYxKJo0plsZqX0kXKSGzzZPRNh85xj299gi628hpgf6b+
E5Cxkycb0gaPZE7audWjLO1444JpYsftU7ij18mhQ6UjXf9CpmXglHHq01+PojeZdd8CeGkXw6TV
tFjX67e2sZdl8aogMCRnjb7xk9kA0KKwdFNhMKh3UBPk7Aa+Og6+zKqfTwPybdS/pr+AF243B/xd
yR2hfOoGylqOw3r5HWTWU7SAkZ4T6ttiw8vUYrQMGD78Vphkqn+UM+7I9n1wE6OOIX3FxQHgKK1a
Py6+a4Lfa7kzJicc3dgcMlizbBhTzJVVDfysZqku4+Kwf73P/sCA/daxHqZGVFMVuNjZXLfNzfVQ
jao0JjotvYrVCTh9y9OGEXeaj632iqDcLG5jVJtgH5tD5M2D8gd06SKMu8h1nMnAV6vCqQESbJdP
EQAErk9IOVoOZPqo2LFNwoWVQrnPoGuTFYwei7ZC0CSJtiqUmGf54lyQgYjHbdiiAB585XS/ayGd
szo4A1b+tPGjR+fL+AYI56kmGHWfeZDpOG3WSVzdxcndG8wFZES8XPNXMnCX4UdwIIJpWfEqa747
X+w0kaoSs9HUFbayC7tuWbc/f4n3WeKNBQktnxg+t5ybjNd4BcRmIobloSLJ7BYJRZhbo+/HowXP
dsIP6PG6GMfCRo2YzS15+g2rQblUehwzHAS2AFTKYQsF4q3guKAfrzzVDeDYPnKC1271ndjBaoi0
ZUedrtGx8ZrNuyA0tyi/fPPKJ9L/9XC4igMwiNXIglapq9aTYan7yAjKoYr3tjojc0tNvlMKj6Rn
3guRhGHTDYv6F7jKKMGlCgjMEVDy/xbxnBP1EW6a/T+k0x1XQXceBMAwJGMrC+H6sCLeemS+rS7I
dAqsRmecxcmj5GQpyw3a11MKVN9kX+U9KblIh+zEvTMe3wNr4imuyw7k8yUax7szrQHC7yzZ17jS
jW7RRD+debdzb3FfpMJaO84rK8EQbg8G6iQPwdfSs1W0f0IV43E71GAYKOxVY/iuhrTKykBqYTQ8
b1qRz9tWvxoweapwctlrcJ0K1hIMm5HP+rT+q1KneNAevnx8xgS/jh5qQbupDB4cBCtHZLc9m1a4
MG3euHT9WppjjvZ++rVxKqCJUoUOMa0Occe7AXgN0MqtnbgB5MqF/Hq7m8K4mywSc9nGZDlkZicp
tTFIdlcnIhBSRVTzL2zXcsos011UtDvd3keUUVgEmuGQ1M16pLvixZ338fygqqdXmiF2fo1AFlEr
YuYp7wakyvhFvBPnRTizFnTCaRykG0/bYTQIQK0aPR4/2OoJshnBj0cyuPgXKOAxsfX5PWyNm1cP
GY+lGK2gzBCUx03f+VOH1oqr1pvXNBitCIcmFRuAGA33l3Y84NRzXtgPE6AFds/zGmk08Snlskjl
tbet1SNZGmMX98uM6psHGnXetSIxv2FQJS9yE/eEuKAB6ru1JRiPjGo2ORii5+bPJk2a1977d5hQ
BZDyNNpcsOn7kBN8BIc52LjQxbusA3UD/iF6AscOKxqGsPo0/z6fv3qaXukiZKquik7DankaUy3K
a8YwtvcnmQ4aKUAwr2uRN03GSOL638z2BJp6up6CEnbUONngZUzNqB4xEjoqiHL5TQDuZVP7e0W+
fq2E5j6o5w8UQmQaQh2bX5LXEXg82i16Vw7iQW/A329XRaoxsIhrAIT5lnkAXiknlgyIhB5r4WqX
RnNej8F5L52obbTwUxmn5qQXlWVGMimz7b9zpoyWwUuwBikVtYdp/dwP+U62O3q2j39VtJu7TzAn
JywCD7fVd/mIF38lBn7s9yMoaxtIuo/20+lK65e7XjD8t+12/4WPMtcI6bn+1IpfLCQD40Utt2Om
W102KRN4jydTqxJ3beqeYLU7UCQN1U4GdH9AEnWePNiUCSaJRKBrdPbeoOC4lV4yYiuXwJ2ahI7U
5w5B6OdoSq97dP4Hh1TmrfE9AZLB3D+qf73adb4YDgiXVqbmQ23qxS9O/+QFom6B0+akzOLNZCS7
K9+CFaJ3XF8Mes4JK9zEONPRmPgdANP5dsg/Gfg883OG6rYgEh/e/9BQ5f5PjLM2WXzM1ruuNv2t
xx1HXolx8pNEW7zgaxlpDop6MpVP56iKWMbdhzn8Fa0E0ew5UPeEYF1+E9265nxzqXZ58k+GQsuo
KQoVT8hN73dHxXtnGHI6hBbsjpAWV7cYwMz26Sga9MnYtSSnYNRhUyNKXjfDFm8rm9bDRBM=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity ps2_fifo is
port(
  Data :  in std_logic_vector(6 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(6 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end ps2_fifo;
architecture beh of ps2_fifo is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
component \~fifo_sc_hs.ps2_fifo\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(6 downto 0);
  Empty: out std_logic;
  Full: out std_logic;
  Q : out std_logic_vector(6 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.ps2_fifo\
port map(
  Clk => Clk,
  Reset => Reset,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(6 downto 0) => Data(6 downto 0),
  Empty => NN,
  Full => Full,
  Q(6 downto 0) => Q(6 downto 0));
  Empty <= NN;
end beh;
