--
--Written by GowinSynthesis
--Tool Version "V1.9.9.02"
--Fri Jun 14 16:07:29 2024

--Source file index table:
--file0 "\C:/working/_Tang_nano/gdp_fpga/VHDL/GDP936X/vhdl/rtl/FPGA/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\C:/working/_Tang_nano/gdp_fpga/VHDL/GDP936X/vhdl/rtl/FPGA/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.9.02_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\C:/Gowin/Gowin_V1.9.9.02_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
h2NufajzsbXKHNozjy19XSs3OC5Pln9e5zhwuNP4iOCH5Xd87cTDinRKHs3rl0Bj6rv8syjk512T
wFCoIsMy4eK/7Eq0s99g+aoacahlknVf/4f7YztAIpiUSSPBoFr2YIlPrtH8DIHFOyI6YPH1LOrq
Ns55/j/iBYHfaX5/fQGZECRSzGSpWywvgBPdFe1YPZrp7z2i9Gn3H1ileKidjd3E1zf+iNl3AUB0
gqZgLtW5SiK3L74uJoUmJPt/oYnA+KFSysYBzHbY2GaiXa+rP0XJpCNzbzzdzLI0DEwhz3ru9HJW
ZF0+7QGS7SeN1qgaj8CFaH2DkqksDnV6snDppA==

`protect encoding=(enctype="base64", line_length=76, bytes=9952)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
omsA5AMwOd1mYdyUo8Slol0qwBpYxFxFEkki9L0tUcvadI6tfQLHHBEXxtwkwUvOSSzN7KRJ0gyh
1/dH4+LbrA/G2ltZWRrGMordIybC8RoW23xHvF4nu8+3v+NjcvX9C7Xgll+Y5FRoNlixuQHcTuZg
LhCQ4LBliLVN+qtLdw8/7RSY5Gsqv1VNZih8TqWdSm1zikxYne6DZrPHmag32rUqi7AWUAL8c0gO
z6TXlJeaXjBvDErtwgJQwykz0rQj7vsqJ0QB1ftKvVuAhhbu2RovfI0EyWHj9ox4vkIKBygVr404
gxlhxtGr/EGDOyMqpnZShjGaarKfmR46j5ax7mRyF3O9Z63vnccYfrTJ9nmmwegDAGu6COllMoQM
Ff16QuFoxyBLGgBZJbIgCFxGBwWCWpyV0aY159/L30Ve3ewwtUS1sHC6ln2Mf4fWwU7YR5vpoypR
qIYCn7va4l1YE7lBNJdiabbrWpCkfikgMytKVIZk57mmcQmbkvhGjSPReASZ6cj6czudXd6KBt1c
oS2zL+AvoySRi16Hbphnb+jR2mWfNjoXr4zM2SZTmvX0K6wrQf02SxaG8XRuyOE5xjbeWntbiMrR
zpWS3sD5XYQkXDGIHpl6H0RvDXeptIfzCZGYrBSZEZFszw+ANLPVLtPbXRmxLKGZC2P2v8UeRWAF
N/iq9+IQcYqETbwlrgDFBV0XVFCebPafo6npxmxGc6G4Du4pae43wHfpn4YwKmmeLRJwF9W76aQc
IdV2nY3JUyakfTzvyXaBFrRAScTEPn7ZmY28Dfs6dxg9oQaSzm0j6HhaZSKFyF4CZtoE8R4Uj4S7
MnQdngd+rGVCtklE+8XVykjRVT/0NDUOvOakk7G9e8lEyCcvsZheQkey/ZZ8/GoN7+9ouJQorwj6
5aaEG8RGi/pMSAhwbcrkRrjHR0Y1yVlOL7PQgSwTqh5/cv6Z9P8+icDUbrnDrSsPxbA0dkfzrtAH
uROFPU9cQH7PecJzItMzzTISo+aeKpDk/tFWq8afLQjR25Zio8tBL7k3leNUzJBCCI0jjpkHzMSm
HKFUXic9j/mqA3fYeYAcXm/Whca3B0Le/oLTVt90tLJIrfVFyzGAubQAZySWpyMOSGkxAySbQeF1
HrmadZxkjVAGCUrAx1XZN8tfA6fHVOruDdbXK7XmxhHoZPHKmN53MQXXptyZUnK6xayVPMk+VNDE
JzabzO7hUIEG2TMi0tX7F5IWnJFOSwk0TF/SfL1ByG2a6yfMdCOpbqkXq8UOvFrlah+TXWhUtjqF
my2YaWv2pwbqKNG3YDsmtu9BAHaoxGPVV2g7BQ2CarFYlrdkyBguFldH4qyGDu2lRhrRNGxt8O9C
Vi9jNfKlt/9z5y88Q5c/3j9wf8B6Cd4IJKgwQx1+MhagoyZf7mu64k7/+0DL0MfABOSisepRFP2Y
B9sNwcD/PIiQxRv/yOqU4TssA+/3anV3mPyV5Tdvxl+suQpjwTOyaiMMhD+U7fTeOTxbITiiz6TE
7in4SSXRFhwh8jN1xyRlnUT/vNEJyp7PTAI4DJarsj3y1docNRZVfcbgjq3lCsZGOvdgMZpyrGcB
BRKae5icQhzq1FCxkbgPW6JOi6ttBTCldy2IZgSQeY2cJJ0wJfaalovlG08dbv2OU3+3yMWRqlTz
PJu3H3igKGUNq3KHpYfcUQykt5b5nqzZUnIhm4v6Qm9BNlBTvIatXp408S2SO49FcjiydxGF1QUd
abjk1Vj+Px8/QvgQOoD4CyXmorVQf0uvQKzRUsV0rCxhJvJAXOXP3/0kH4OO/aXuB469yjH9Po/h
h/0N16rVu75VtQq3wJKkJA1lOdqIkK0gUGSVkw5swYcQzb/PcPLrs3tetQpq5g1hCoDOE/JRlfC7
FkkxDSZrmN60tWKe5OYhClFOociM1HFL49DDVsybYk1rfXYdjalEfnp5k1nq7aMRBU/fCp4o+vBm
DKjsASGCTph+YGbmNdh61WPL6Gr8ftYrKnKY7EhOI8tFI3dMBAzRGTCk6ExVsS3wRK7GvStXjyz+
016df7Rp0jn51Lwcdhvm6SBemCQzLVnqJ4OJgz7zuEzWq4NBZ5XbEO0MG5z5EUv9hF9mA0l5iGAt
pQdisrSynrJFAt77qhlncfrwV9LIT57xRobSqkkRk79+j4CvmOQ9sWn/ZwvIixKTGQWjXs9QYScr
QQF7O+1Q0x4A1PTG81ZTGCbDYV6Agsfj00/YWHLo/5mjBsz0W76yTzVXu3vvfwGiKK0ZXIfwrt7W
VZE+1fCoGL2LlDfFFT+EF549A8FcB4LjNnveQjJtm2OgX89Bv1dqK/B2yj7CxIwrsfNBEmjRkEjh
VoSu5X7jZMiLCfygz4En6lnKQxPdFkbAKQ3ZEdnr52cnRxr5SnJ5J8r/Kz4KxuVMaF594HZtWq9F
k2Axeh+xR+rtW2Q/VD3hBG1dRXQYpQ9rCad5hUr9X9I3uuoG3ssWMS1ObDN+I52KDFUnskchgtbx
kcDpPE0SHZqjnQOf2gsa3cZ7L7UF+fvB7WuQoMiMrqfhJ9VcU1jqbB+sLEUJSZIO3kkgXu99S5bR
eG10VQ/miDZMXDM8TkJw4WHiFvU+lddYDx/18lYdjP6a6CLbWu/VjXxRxgG/TQ06l9FEvHcdixAd
YuPVXFvmpI3SmEWawT/mZyydoMBSrYthxlFoNn3KiA4E4TmB6j/hQ4hs1QzrhPI6TYzk6/6iLpvN
FIDUeP6nbPbOTCUy2UDvD6CcDpVWOIzciG406jBhR0DyyqEcadd0hjN2Fd4t+uJu2evCtFdNYiLQ
H2yRwXZY4hbFi0bi5NEtu4LubD5NqYtiBZFFeN4DRn2636aC0HRcQfUJHJxdlKU9e8wf1PqjJYrE
FFppe9jZaN5IzuvKOXk+/e/a7+LbXU3R0jyYpVbQ34Mkws57g52ZelfuWv6QYP1kHsClys0c74hp
5k9BVWzLrJuWBMe/n1GdbOQCX05Q06vZioDULeA0GXvycSf6z0uGU4l2Yn8DcnA5P+yMwSag4YA/
mOug68j6b42LvjfrsI/lWlfk7/G81p7upVs6UbwWNhVCZJ11woK5NdfTPfExNTvCZsblqz+6mltl
3N/u74AOPkg93m4Agt1YRL7gfLhshX2ojfl99mj4ZHdS2xgG4Bn+fgr4DRirOM4hzBL6b4mss0/g
Vzw1WjevKt8At/KTIiCgID3ksY+zV6M+obbGe3heHiPCM9qqYxd/dAYDQHQGB2F4huZLDbSuqR7O
zMmYqZ0lDZ1dTJqVTb3PmLE6etKZJuqGcIyuFmKnKXYbjQZLY+dmciEQ5ahYQ83tgUxxNljWvSGc
6UxUY8jL9uMm3kcoWyfo6Tp6u3cyrjAJ7fUgZSUzzpdMAKEHEIb/oXLANQGLfp6TWIMSkpskSpdM
ASCSJNMbLC4yYNYA17mJnGti7bstia73CDUBgyJl32jRYa7XWgsLdGLYt1g7zvYpTaHwYXd5tzn5
6jyMs8jrTsKLDnnCfbopb/fxD4j04s/p6YTo4TgZEGX+AsbF7mOW+4Psn3cgt9yfBXseXXlpe4L5
4tkrthMDii87ExfpQb4MqnebCV/QSEvvvwGzMeJ8C4SWX4X1tPHaLWop5Lgaj5+TfbSCdXnal+nY
DX3HAmQ0bVS0rDVf2pI61yvli4F2o2jvtlBQFCv3ox7HKgMIe6/E4lqD7gnnBO+rM0lJ+YQIGbH3
egk69z0yZ7nXmtOzPtGb5ukOYN8HR0UiHkjSXPNwYXUtbW1axYbMlv7L8QIZb0kamvabVhTaVDAq
AkPHEjOFJgVOu2yQ7OO8jVbuPpCg42UO5C2UI60cjevjnaWSXepqhG+m39I59BrCinQ4F2sdhqRh
NBq1zPpWqE0kwH2NmYwpOl7tdrzLkCPWq11MNvBGkRo0mdY3UrEFEmoseQSX6ODcMc0pPH7IXC/k
jP/OGpF5fu88sUV9QyImooNZdWhumvoBKidXczN+UJ96lWvV6isJhNlHzcgUes1BhFadxhfXRGFa
Hux+fhemFlgPvO2i7YJTyB9eMQ1KWRoCGqYRgdCBXtlgvtfZFiTH1IezGGrsKwdHQYEd1TMr9JG6
i1u7/5z67cp8zkD2yfGXo0QemGvR4sLbtgt5zZWysD0y2Vz7TIOadEhUWT7O5nz4F+MkGHLbkjui
q8z57HAcVdsBxnDoUQjJFxKuykPpG+qDm9kdzEUmBthmF0zlPQCF2usPdlSEwzThxmVdSU8Ieupv
O1p8UAxgi7WFiOpm+ft6+TIEFR0ntTrdSwnDO8hM5gfuAy6ZXiwV2MgcqOUgUIdfglxVKQZvm1os
v5DysZKJMSU6t1eCEzbzPWL1lvzrapajFv6fg5PgirAriGCJjv38gtNNd9ecmKNqqxjCTsy9r59n
cm+WMga9uSqCjr4gVeT4MFwkwhbUa22+/cdlyGZfy83f10WE1ztyBuoJs4b2RtO82bdgJ1j/8SZZ
hQmUALInhMciq3E0jaMMfnEaQaaTd53yFS6gHFX2zzDA7KAxZ6L8iYMjFw19UkKD46uRmGQy1GSL
8MgnlQufnYZ1/Uwmq6I7xtnqj4/4KSZu/lK+TJXMHoANS0ZyJSwQ2vtL0gL3MNsyhw7olwaJNZMB
dG5fr9be17svP7a6W0UPAyW0+lRmAPw5eLMBsiC1HnL8oecw58Ye/sP6uWRKwQXfZ7FttyRe5uIy
rBdESffQtanBFidDTxSkcgB7Ev/g0zKxPoMGEV7/Ab058OTErEsAv04NfGgbz0uxrXXUsnmt9A9h
yMPBr7L2lYpIFNQjSMVJHMAiTOlqtGncez/B2JU9XhVjRGsfS2fRE7nEtiRdaY1WjbkVCrQi2F3h
hLyqLGeLgzcE4p+7N6pAbSZ/KIlNMax3C07FgAnnyLgnXUmvG0QP3srm2WwxLfV7zGRnLFsvFVPY
VLWL8Pr/qYOxKVoZDOvrAm2XOjnHyvyAQnURgSb7eo2hTiinrd92L7Vesl5NwxJE3kwmcHJQdHj2
Yniwlwm0xKyITuGY9tLcOsJ59HbSQiLwDiZzGi3ZpehNYiSKciVDhnyYPGdwSJOtJguKfklbrk+q
0OQF1kNE4OAkH9wxE+0GsIT9x9J4yM2BSj7TzGqGOTsi+UB/GtceYzABC0jBFCK14eurx7+MR7BA
Ky3bNlGZv/+75PDjGsPfQ3i+nKvao3RxGPjMhCJOCN1mRBPAXW/t7C0pTNkG9ck1yXXM0TWGdBjY
Jqk7eSWv/BpRdqi3+0MGa5SwBMeobOQjHXOU/nhJgPyetwajVz5pmVt8UABb6551s7nP+T550Hya
oG2YLaaEw/JU7gx5BOVHl2UIDt7Yrh+C9w0hEb6I8FXLu5ySnT7a4dfWCgsJ6agvevoKbuVhWME6
YyhTFt3mkpRU+mghuZmgBviwVUpKYm6cKkEutAMm8jrPtn/rPufP8DpB3W+UZo4KOGWRHCmKhNYD
Yen3H6xU9OjrmQUCVTPa2OsZ4Smi6tEPT0yO+S79XGo3Vpj4r78HsVXKLp2tuDXp3VAE4YNLaZ2j
kTEwlZPJiKWvnGrAUFOvo7X94IpF2WLJMWJk/XwYWNdekoOcDyMcbmiGhNYn1KoI3F671b7JBhuS
7IfLqnXzZreKhHGMZcfjiOwwTskF28O5W8UmMgOhE7CZkZQHkh9FwqtUI/BFHIAy5sBHvGhTEIgf
2W9nPsI/tvccj5bGlSHDGX4GX0lJYUu9x5brLylIpT2r11OzxxFaMym8Z/5mi3uOYwLvTwySt3RT
uCpo/aTjLAFHOWT4k6+l+Ji3Im5slVHWhJouwoKpfg0KagUE2rywe8ljh1AEu7hNZ4ZRS6uaaFjG
3y0LEKCb0k3HNpA96yPMAGlckUhoU97UH3D0G6MlKTmM2ar6lKbYnCCdwbXbscP/2aXDys/2H/Yx
LVWMzCCItt2U7wR01D46dD707ObiY70Sr25K1WzEMWxfUHG4ksMWGz9h4QAazHDbpkL6miXwqNfm
UTHWroTCAxnTxfIs4Ld5l9CrwuugSMgJxitFeUK1eMTJgU0x1QxGL1K6VGc5ucBEz8iFY4WyDgUf
np9xuo3mHZq4nJjZ8xiqMlMEKJrlR1aztvzracDP8JrDuPWN+NeyGf02MBuc4pogb0AK6xjPH/5T
MnyCYx1SczNJU4iY//4cRLrXOK6xv7RU/ccZl7mIl29+hT2zchcc8gsd9znjmrvAfkCO1o7mfBKY
cZ1P/coqoNoDV97KqlSa0qleoTlQmiWOD88+L5P0Py90/UsCNtuMEIM1v9utH6jQrkivEArWxbVp
qMdm4nEaGOTFH2ul53o0bW/vUalB/qq4mdnfVMIAWBfeiL0FWuWDHi/VuL7ysNHtwmWzLV9a1Y35
kd47byGy1J4PmzNZFj3Brm5Za+TqUHhHVGZQOhCUoK8csXLo18swxkZApMwPoPqytmu0+NlO8fyr
k38DZjWySgdSpnCIh/JkSW7j/x2b9n2Igo+/WHjU6Sc0+TIeOzESjx/EACgijkz2xlxWd5ZS3uTN
PGA2OH1V7tkckfWFs+HzqlT4a0AXAYIYd97pH40QRbprCBron9dekzBclIcgcLelIfzDkRDFTvb1
xbuQ+ndxdmH/6myv/uQdiN6kdM7slH7Aa8i4zt/MuoIsmZtu0/Ble/6ycMs14LOwsu1QE3XQCp64
FzQ1AT0JEVa6Nwf5px1WAARGU2zldEEv8V49KiTzdmxDuzoRS87X9W+R/hbsWIbhkSb85nkO1a4D
/E7/yUWiBvxKfYK+2e/Q04xb3Qzp1pMNWm9607EW7mCiz5IDglaCfMsvq/n/5RtilN9pJzhfEIQS
JllEYYZCmpEeCSnTsDeSGYEJa3f8EhKaCW4jcOvaNwU8cwd5Y3/9np4op3+JkWYO8Wjv4P7LIcgK
J/Z8lo2hxU/oOoa3pT50jOKoDM8YX10x0PDXD779eI3ABxdaW/CjGFaCn9OXgQAoNbNDIeAYdEoy
uhbZ1zEpzp+CBGURc3qVldkulXyq/Qa8LFROB/0n2yvVmWy28tgsJpkVedSIIBeiNGk5Gppj4xmp
LFSszNhlJnvShKMHEVcVbV9Fwve8nIkvMa8Qa2uctIYdzE9eAr3meIh86D4sM/+9v0KUjqBA0wN6
XZPPm9fiyha8tnP35Y9WIr1kJo8bthJ0NZfVa12y5gXkd+FWeYDgV1lfcZXfb2W/qbt3P4JmVgkA
MXVCXpoj4DBrdR6ldmCADWRFof8hlOXdnXpTQkZ0M5+Gs1Iy+b+cUFVCwpwn0b/ppCQ3wqWTJppB
aClaqPds6fzexa+xlnDqVh8aTszW8pVL3PpGFWVi8BCPZ7yr4vbALcB6Uywp/FjOcUt+u6Ez+K2n
/8bNsOk9oNzZCNcJDaduc/04YOt56VJUYteZ2FnHzpKREPKnJ/eHDLMD9Z7EIMAMxhcfZhLk9Ylg
8I3tXiZJRULgWfq8JACDqAzfBPbdrrk8lA0E3KbGa1KdTaRJO7jlVIbA2ark6SK8v3jCwQwkvQm6
pvlKQn0CkCR2nW8FRKguPGDqlXIlJj5YeLdVpr6F2HqYGailh01LH7yKlQwqptLbh7F3jjLYShu9
SSqhVk1mEW8xip60VQhQAwk8OffcWMF9h4Aqg6bgKPmrY+7YqXIN6lrVPkd271UL+Jli9MciUjkx
ly0tXtzNICCZHPjzk6OEkw4ZwdjwcgkhSz6afRJMWJssPBFvG7f0nrxa8bZqr69O1n82iW8uNtFX
5EB+O+dKImrW6Djoy0XIYd8Q8jqhmNbNexxX3idgfDZtIpjusL29pg5Nau6y0+RXz7KtHw9nYCZl
diw1GPeKANs8dGZl+Th6gJlHBgoKQWAx/Im/hvYBYgBNBaLnqgDgSXXw/LdAJaiTPFUXX9bTe2Lc
HPpWjoKLzJlilufo9zz7cYaX1sJ6oTZ2wwSS+6//McEHUvG5ONT+Bm6uxbU4v8H+Wf75/x3fMWDT
D6Dz4VaoRujZ4HJTDVdTR0XXS5qOsXgimCu1w3bK7IH7qJ4WNbNpooSYH6hTL+ve6he6RfTGXvO7
9fwONec31G47vWdJbsEZiccPTaQjzBekY6GvCslqZWDWlkM722yg43Pu/jcUu4aGd/rM2pOeAsS6
yQBpGD79WMtLZf7hZQhPl4yQLIMF8hb9dcRUKqcA2IKXcnojczRcN0V34SFJohBW9GAbL8/JKNym
yRDrRDXN6l+6E7tceEo4qZMOW3385gF70i/GldknWg5SguS5idjZ9KcOzo8IAY3DLafd5m8nQCBA
gGFLyZZvAORPBj6zu7wqAhOBu0hjpqxt6k4MCHyOfT89ueWdRpRddCCVk6hC9arUxv4Ths6dWdSv
cW5p59MaWSxJChK+3x/j4quBC8UF9va7vc4oUyqwpHk147xCZGbXli8dOo1R//xq+X1RB2f+WDCf
5l7iWuEP2aXVya/pjOXKDvSIJBlXHiX2PndmiiujMoQsBS0iwwzIqBlw/J30yFAnrV0kKaagefe0
5NvlswrlkU95ceAENsmjYsyHFQh1W/OQLQPKXoLBoK7bXrYz/qMTQxcCq8SQYe4gJAJU6qJMltKk
KDCgeA7diZjM+B81gHltdanmug2MR7LIMd/BG3Nbo4d6E6oYnaN2VqYdy/IiXue43kGBaE/3pn11
YX2hQjqhrH0kr8cRFdglmf07+apzunEr2dWoUeloElfKlELB6c4MqdWXvZIUg6zhuZObuvLYqPg4
DQIXUIgOS9G29md2+9wX1DX+mHGWwaYleR7VbO6gV1gQbfT7sTiIHC7AQi8esNOhOfgDHGdMCRvK
ybWX9J0Q5qgmeiK9uSAAoc+m/EU7OE7SRa28iBo4V3Pew7Nj75TSa3BHhfFOYwYlyggFZa4N+pt5
KuAlg219UidTYQAuQwXxi3KDp/wCPrDAeHFwFc6IBbBIURQlRpNn7N+o4aGTkEMzBuBX06jyR60V
l9re8XMrZ0ZIIoyOa/pPt5NZNOhxxVeTs7e7cLJ6H9Jv9Y67/tEmmhABDVoJF64/omikeBJeB6pT
tlHv2n5yLVG8TVZ261/oEwvGpr/Uznvjad15sffS33W9A4svhKrlSz4MENPAN+37xTTdg2gMWawZ
BTnFKWNkdO1gTHLvUcj2IPmLEI5xyADGJZ+54H0NVJ5cWv3U8fvrBglvd+TFccWvuQ4horWiSgbw
TH4dDwPXTF9SaHEQPyR5Efn80wQxg4AIe4yLH0EcGIjpprF8CC7xHHw1fdZP+ieA9Js98Zz8Xbc+
LxeWplnHM/mwq6BDKHWteWoMOSLOxQRw07BF558b0NFzmyRKU1ZDVTniyhmgLmqlxtNdJe/Zrelf
ZvsUbTAbehniefhGmXwFy3faWCcUSI3iVurkFMZaZhI/pr79zH/EoryBY5u751Lf0/c352cn/Awx
qU2AdVQn9+ZVEYq4mYdD5npC3884GfOdotS4e73sn2SNsR5NyRDNCnIU9b8j9itHMOqY8CO+c+l3
2WZqu5eZX86n3IQEpYAjDWH0YNO6k9/s5g4RvqnuT8AsWWY4fr1pA/fDM6BWeE3hucWY00601KEI
BPasSnKpaBCriwVvoV4Eg8YMr06zOmSzzfu6Qt58FZ0TsTZwQkBRebZi/xHqkgimirvZYkt24HVX
5707WFFEr+ucaT3eHvjk0ElDcmWEh9sQqCC/vteo86WStzVK9uODRD1AtFX+P/CcEOUZ4GVhmLXc
2bKhrtvSurH8EstUBxOTtuav0cc99MQv7SN6ZkWxNRjPvApFrT+5L8LXdlLalmJQymh8XygREAO/
qQB5dtJ5lFjv1KVzw0/REsDWWSg3r3XwZwWDzKflT9wJfJ6e20GIDHIPtZ3Cm+z6LSxxOfHgEk5c
tWFs0z03pl0YC+ZTofo0LR+I6tfv2jhVA0hCLpyYvJbSHy+V6ppTImR0OwBWPLch6L8TvNrRWjcK
GR+WHiA7sJepvVDoZgzWsy0OmxBB+UMtANzc/Wz5emIzCVcAIh/hzykDXjmYgyoHOgAg2rvMEMqo
TBAyrW1G2A6swsmcGooKIRkXBoQkKF0/8T3RYsDJq7kO4U2u9o5VFtxRdGJ+EJvtSCMfHen/YQy9
VR7tcODcGShJ6jmTfX3ZNbFC/XRYguqGbSfIv62D9+80tyIOIcxz40Sev3KeqhqNDkrC1Scmt1Le
QyLx4HnnfKVbK7BHY75IwGHDU2LrjQXAAjXX/oBl90+qapWCMOqkHcG4Kxt+alUcy4pqHKypBX5f
zfDX4OgPcSkCRO0EFbQgsWnAonlDgYYgcRtObdyAOvxTYqWRNry4aHoUo7WBBY81FyQh/AqkmRb8
ikBY8ughVjO4xJSSpCON3/9OwYCW2kmHa6L25MSg1bplt3IEifgZjUDGODT/uEkwxoY2z+AU+sLU
1vT0HX0Hg4IsdW0iH2/M4n6C1Gra4O7kr7LPEz8qYiOuWM8KeKLN0JbdDs+NYtfSEpexWS6Kpaqy
/aNgFbaPKynysSTylKT8TuPkw7TZo9NpRM/Io/G4we1kREnY1jizlV4n4vKgRFhiIfW+Z9oRi52V
W23mWEyoqek8cobqZOat2Cnr2aCb3n5k4FEI3cwvv2PgK/aMgcoz7yO4HM66A+uBuGX+G+oBiVBJ
PQi4vy77DiR9z3ytWf9mUPiJaPAFuzfEnceE9CNX/DyVw9AVzSG+Pc0MyvWeEsrkOlZaySxsp301
/IbqeQlnlrRIR87Imwul6xmmyaBpY/M5Jm3+kZmQJUt/temJXNgxv3s47Iu4LZvoWWXj0w0fNwCi
sqyOY2NkZvXGak2F0Uf7p+/oxa9faLRaviQ5/PgLA+5+1GG1K0/6EIO3vsYsSqF6q2HtCPDGnxoP
5amu9Q9iyvTuMVhgjGC927HZ0NIJEuLY4lWY0qUmCh5bLV8tkI4MTAVIK8p8HpPU+Gd6NTo7jAL+
CKwSoPSBEE2PbbMJ09heLUU2hYQy4Dv0n9gaApxBHYSV9eNrgSUc3Aqmo/ehi1zde6w6Wrd+dPq9
I6dW9FOPQmu9XewstyFZgTS+g6gkdYWr0O8hbZqQok3XtPWM2Z0jxRtKYjU/1az4Y8mK/e4fdqNM
vIjhk5GSEeUHnNMch19fwgi5xW613eW9RwLhxKYGiTPFTSRoTbRFlwaSUZxPGnu9f2ihcGJTWZU+
J1WJL7K5ujklApTaP9RmbEX1zGnmXhLujrfVUSz0f+qDs276odXWvS+dusiawhfD45OnBoIwqqj0
CzKNEOLfZWa5AaEHymDaVZyunxLAaJHkN2ByrE5qvhyBJ7ZeW60+am+HPBnJs73C4CWFzkVr9j19
Yv+sFu3tDV5MihYwUTkoMYv21pqfNvFO265M3pwctj/kyRz+CZ81+II/q9JWLKjjd6Sq9yqFtFZr
EAsC9ndO2oGQ99PetLapTBtYSDJrjOiEF02reqZn6QzCOJzpbXCc/X39LkjL1W81VXFRXpjBzbrp
KRo32Jh7iT7RIfV6Py7lrWH8/jneMl4r8iLQ1fNXRRWP28PvS13KBrw7br6s1g8wJkQ+/s+ZXc5s
GNNJ3kvU0RGgBL4Qxgsj88bqxdBjzedevFE8dDmGlQvztyFBSRnUCpoBcHWQP/UORMGGO2Jo0kfr
lWCwUAFGMozFyyvhKnc1zVpGucDaAp9vrgpphm/QJBSIoXYkTrnMFlc5q5nNxLI9KSlPR9TAbD0Q
bXeG9MA5DqxDQPmEEo/cL/jt54mr2lGFX6ZJbwZIUrVZCuLa2fqNvSTxcAeBE6dlt0w++MLuxJlB
z4DQv9CR/5s/RGN49qQFJ7MR5PH7SGl0RjlQA6hrTKLuCvNChdoYhHEjbDM/Z+TzlqyywOF/Sixb
iHZBJEeN0mCMLvOMV6uV52rz4YeZ2Mbb3ush3Of8nzys6bDsUUpG4Q55RMQM7xbwmL4fcQw+jUu/
5izsBjf7ba5sUXode5gFLkpN0Qy8dhsS0j6fQg/toC996aWYr6PfjlNPahemttZkTOhleTcXV0EG
mW80dBGJuQ2dKykS2tcistokhC3J9vdXwP7m8tK95PWFvcx3uNkGwaMy1oBD88MxexInxCurvAEC
nJ29hcuSm0S2ItMYiPLCjSwgy9XD97aBzUtnYs0+grORNZw6r1W2IjmNPQxx411sljdi7hKrYOEg
eSKkNrmW0Exj3OBz3gP4SeMlXWDbYSBrGC34b1KBWoM8sJnjAevV9CsZBdub5eLx991xsZe+VOnp
uEn3FgkeH81Nb8XbYb4DV9HL2IdjcUCPa0TUkDZAwbvfjCkmwu0bl8GjGFDRcsCK8f0h+uMd5bBJ
IvWKv3cp2VJdvsMDCVQ5BDQ59AyAIbNSjtN+vnChea62+hRoDonvCrMw1EhGlZwmdEhVEJFO2wNf
8By+ke2PV7h9HhKLCDVEZln4cGRCkEi3RPFB32m5EtSsnephYHBcXEppZB0z7aMzZCr/KE+p4L9j
EynaaudoPipneviSyxmLGSKbNkpsriAlTUWGJHBBc69bJF60D9zLVXHMamDFFzQZDk6DpLR+lWX7
v7hzJmTGZc9RbC13cfOKsUYCsiIFmA+ZkM93rIIIugyfqSik2OIF8sU8w7B2daNHFcn232NIzkvU
S7nNxC8vTGP9Va0ab4J93j0V5bC6yT2nbrp2DGlQq69YEul2MBEdv7tA7OX0Lu0jXHPrblLMFjNG
Ggdo5TxtdELyAcIYh1jWaO54B5Slv8o45BPJ8g2SA0XBV2HLOYHditnNodcCzX678YWSyZ28tnuk
qUjbP8/PDcuIVGkcmDJP9vzrmZ35viUkfyUAo/vWSuGlZdDpYQcDhBfcYALF41JCtTsR95whhZJc
S7hOLpTymrZhBP1lGFxN2+xJrdNvgEU/4XmbyVehiVt2FPGfGU1VlDFdAykdopPZrFtw90tqVz0h
BH6Ljsj5sh6bHLX7OkQ0muVkyfskD2nNh+5QZ7KMGjuAVSSgKeXwwvqHZpsHQNXpS5vFQO87b73D
Z9IUB2DwuMGjecu+Mhb9xm3IAqecms9Ns3++NjiPra2+7vTdJ1SOWx0m4frgD/h88jfZY2NJyI/P
KinLQv0roaS1W+JBMvdoAgXTn++c5hc6ElLxK4P1NR/s/1N1+H/VHlJJLCEVE9f5S7uY9FoRpmYf
k+Fdwn7JHbiEenfoDdmSDVWUTllPenvuBf08FBcFbrWBpE4k/Z+P0qUk5yTwPJdyMxXolArXduZN
cxHhkDg1v6IbU1SRIbAjWeSESbtEKR54xAAOweblikuy/Q==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity video_fifo is
port(
  Data :  in std_logic_vector(31 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  AlmostEmptyTh :  in std_logic_vector(3 downto 0);
  Almost_Empty :  out std_logic;
  Q :  out std_logic_vector(31 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end video_fifo;
architecture beh of video_fifo is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
component \~fifo_sc_hs.video_fifo\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  AlmostEmptyTh : in std_logic_vector(3 downto 0);
  Data : in std_logic_vector(31 downto 0);
  Empty: out std_logic;
  Full: out std_logic;
  Almost_Empty: out std_logic;
  Q : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.video_fifo\
port map(
  Clk => Clk,
  Reset => Reset,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  WrEn => WrEn,
  RdEn => RdEn,
  AlmostEmptyTh(3 downto 0) => AlmostEmptyTh(3 downto 0),
  Data(31 downto 0) => Data(31 downto 0),
  Empty => NN,
  Full => Full,
  Almost_Empty => Almost_Empty,
  Q(31 downto 0) => Q(31 downto 0));
  Empty <= NN;
end beh;
