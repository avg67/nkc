--------------------------------------------------------------------------------
-- Project     : Single Chip NDR Computer
-- Module      : GDP 936X Display processor - Color Lookup Table
-- File        : GDP_clut.vhd
-- Description :
--------------------------------------------------------------------------------
-- Author       : Andreas Voggeneder
-- Organisation : FH-Hagenberg
-- Department   : Hardware/Software Systems Engineering
-- Language     : VHDL'87
--------------------------------------------------------------------------------
-- Copyright (c) 2007 by Andreas Voggeneder
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.DffGlobal.all;
use work.gdp_global.all;

entity gdp_clut_256_24 is
  port (
      reset_n_i    : in  std_ulogic;
      clk_i        : in  std_ulogic; 
      clk_en_i     : in  std_ulogic;
      WrAddress_i  : in  std_ulogic_vector(7 downto 0); 
      Data_i       : in  std_ulogic_vector(23 downto 0); 
      WE_i         : in  std_ulogic; 
      RdAddress1_i : in  std_ulogic_vector(7 downto 0); 
      Data1_o      : out std_ulogic_vector(23 downto 0);
      RdAddress2_i : in  std_ulogic_vector(7 downto 0); 
      Data2_o      : out std_ulogic_vector(23 downto 0)
   );
end gdp_clut_256_24;

architecture rtl of gdp_clut_256_24 is
  type CLUT_ARRAY_t is array(0 to 255) of std_ulogic_vector(23 downto 0);
  function reset_f return CLUT_ARRAY_t is
  begin
    -- 256 color ANSI palette rg. https://www.hackitu.de/termcolor256/
    -- Only colors 0 - 15 are different, and there are only 6 grey colors available
    return ("000000000000000000000000",   -- 0  Schwarz       
            "111111111111111111111111",   -- 1  Weiß          
            "111111111111111100000000",   -- 2  Gelb          
            "000000001111111100000000",   -- 3  Grün          
            "111111110000000000000000",   -- 4  Rot           
            "000000000000000011111111",   -- 5  Blau          
            "100000000000000011111111",   -- 6  Violett       
            "000000001111111111111111",   -- 7  Zyan          
            "010000000100000001000000",   -- 8  Dunkelgrau    
            "100000001000000010000000",   -- 9  Hellgrau      
            "011000000110000000000000",   -- 10 Dunkelgelb    
            "000000000110000000000000",   -- 11 Dunkelgrün    
            "011000000000000000000000",   -- 12 Dunkelrot     
            "000000000000000001100000",   -- 13 Dunkelblau    
            "011000000000000001100000",   -- 14 Violett dunkel
            "000000000110000001100000",   -- 15 Zyan dunkel   
            "001101110011011100110111",
            "001101110011011101011111",
            "001101110011011110000111",
            "001101110011011110101111",
            "001101110011011111010111",
            "001101110011011111111111",
            "001101110101111100110111",
            "001101110101111101011111",
            "001101110101111110000111",
            "001101110101111110101111",
            "001101110101111111010111",
            "001101110101111111111111",
            "001101111000011100110111",
            "001101111000011101011111",
            "001101111000011110000111",
            "001101111000011110101111",
            "001101111000011111010111",
            "001101111000011111111111",
            "001101111010111100110111",
            "001101111010111101011111",
            "001101111010111110000111",
            "001101111010111110101111",
            "001101111010111111010111",
            "001101111010111111111111",
            "001101111101011100110111",
            "001101111101011101011111",
            "001101111101011110000111",
            "001101111101011110101111",
            "001101111101011111010111",
            "001101111101011111111111",
            "001101111111111100110111",
            "001101111111111101011111",
            "001101111111111110000111",
            "001101111111111110101111",
            "001101111111111111010111",
            "001101111111111111111111",
            "010111110011011100110111",
            "010111110011011101011111",
            "010111110011011110000111",
            "010111110011011110101111",
            "010111110011011111010111",
            "010111110011011111111111",
            "010111110101111100110111",
            "010111110101111101011111",
            "010111110101111110000111",
            "010111110101111110101111",
            "010111110101111111010111",
            "010111110101111111111111",
            "010111111000011100110111",
            "010111111000011101011111",
            "010111111000011110000111",
            "010111111000011110101111",
            "010111111000011111010111",
            "010111111000011111111111",
            "010111111010111100110111",
            "010111111010111101011111",
            "010111111010111110000111",
            "010111111010111110101111",
            "010111111010111111010111",
            "010111111010111111111111",
            "010111111101011100110111",
            "010111111101011101011111",
            "010111111101011110000111",
            "010111111101011110101111",
            "010111111101011111010111",
            "010111111101011111111111",
            "010111111111111100110111",
            "010111111111111101011111",
            "010111111111111110000111",
            "010111111111111110101111",
            "010111111111111111010111",
            "010111111111111111111111",
            "100001110011011100110111",
            "100001110011011101011111",
            "100001110011011110000111",
            "100001110011011110101111",
            "100001110011011111010111",
            "100001110011011111111111",
            "100001110101111100110111",
            "100001110101111101011111",
            "100001110101111110000111",
            "100001110101111110101111",
            "100001110101111111010111",
            "100001110101111111111111",
            "100001111000011100110111",
            "100001111000011101011111",
            "100001111000011110000111",
            "100001111000011110101111",
            "100001111000011111010111",
            "100001111000011111111111",
            "100001111010111100110111",
            "100001111010111101011111",
            "100001111010111110000111",
            "100001111010111110101111",
            "100001111010111111010111",
            "100001111010111111111111",
            "100001111101011100110111",
            "100001111101011101011111",
            "100001111101011110000111",
            "100001111101011110101111",
            "100001111101011111010111",
            "100001111101011111111111",
            "100001111111111100110111",
            "100001111111111101011111",
            "100001111111111110000111",
            "100001111111111110101111",
            "100001111111111111010111",
            "100001111111111111111111",
            "101011110011011100110111",
            "101011110011011101011111",
            "101011110011011110000111",
            "101011110011011110101111",
            "101011110011011111010111",
            "101011110011011111111111",
            "101011110101111100110111",
            "101011110101111101011111",
            "101011110101111110000111",
            "101011110101111110101111",
            "101011110101111111010111",
            "101011110101111111111111",
            "101011111000011100110111",
            "101011111000011101011111",
            "101011111000011110000111",
            "101011111000011110101111",
            "101011111000011111010111",
            "101011111000011111111111",
            "101011111010111100110111",
            "101011111010111101011111",
            "101011111010111110000111",
            "101011111010111110101111",
            "101011111010111111010111",
            "101011111010111111111111",
            "101011111101011100110111",
            "101011111101011101011111",
            "101011111101011110000111",
            "101011111101011110101111",
            "101011111101011111010111",
            "101011111101011111111111",
            "101011111111111100110111",
            "101011111111111101011111",
            "101011111111111110000111",
            "101011111111111110101111",
            "101011111111111111010111",
            "101011111111111111111111",
            "110101110011011100110111",
            "110101110011011101011111",
            "110101110011011110000111",
            "110101110011011110101111",
            "110101110011011111010111",
            "110101110011011111111111",
            "110101110101111100110111",
            "110101110101111101011111",
            "110101110101111110000111",
            "110101110101111110101111",
            "110101110101111111010111",
            "110101110101111111111111",
            "110101111000011100110111",
            "110101111000011101011111",
            "110101111000011110000111",
            "110101111000011110101111",
            "110101111000011111010111",
            "110101111000011111111111",
            "110101111010111100110111",
            "110101111010111101011111",
            "110101111010111110000111",
            "110101111010111110101111",
            "110101111010111111010111",
            "110101111010111111111111",
            "110101111101011100110111",
            "110101111101011101011111",
            "110101111101011110000111",
            "110101111101011110101111",
            "110101111101011111010111",
            "110101111101011111111111",
            "110101111111111100110111",
            "110101111111111101011111",
            "110101111111111110000111",
            "110101111111111110101111",
            "110101111111111111010111",
            "110101111111111111111111",
            "111111110011011100110111",
            "111111110011011101011111",
            "111111110011011110000111",
            "111111110011011110101111",
            "111111110011011111010111",
            "111111110011011111111111",
            "111111110101111100110111",
            "111111110101111101011111",
            "111111110101111110000111",
            "111111110101111110101111",
            "111111110101111111010111",
            "111111110101111111111111",
            "111111111000011100110111",
            "111111111000011101011111",
            "111111111000011110000111",
            "111111111000011110101111",
            "111111111000011111010111",
            "111111111000011111111111",
            "111111111010111100110111",
            "111111111010111101011111",
            "111111111010111110000111",
            "111111111010111110101111",
            "111111111010111111010111",
            "111111111010111111111111",
            "111111111101011100110111",
            "111111111101011101011111",
            "111111111101011110000111",
            "111111111101011110101111",
            "111111111101011111010111",
            "111111111101011111111111",
            "111111111111111100110111",
            "111111111111111101011111",
            "111111111111111110000111",
            "111111111111111110101111",
            "111111111111111111010111",
            "111111111111111111111111",
            "000010000000100000001000",
            "000100100001001000010010",
            "000111000001110000011100",
            "001001100010011000100110",
            "001100000011000000110000",
            "001110100011101000111010",
            "010001000100010001000100",
            "010011100100111001001110",
            "010110000101100001011000",
            "011000100110001001100010",
            "011011000110110001101100",
            "011101100111011001110110",
            "100000001000000010000000",
            "100010101000101010001010",
            "100101001001010010010100",
            "100111101001111010011110",
            "101010001010100010101000",
            "101100101011001010110010",
            "101111001011110010111100",
            "110001101100011011000110",
            "110100001101000011010000",
            "110110101101101011011010",
            "111001001110010011100100",
            "111011101110111011101110"
         );
  end;
  signal clut     : CLUT_ARRAY_t:= reset_f;
  signal Data2_s  : std_ulogic_vector(23 downto 0);

begin
--  process (reset_n_i,clk_i)
--	begin
--  	if reset_n_i = ResetActive_c then
--      clut <= reset_f;
--		elsif clk_i'event and clk_i = '1' then
--		  if clk_en_i = '1' then
--  			if WE_i = '1' then
--  				clut(to_integer(unsigned(WrAddress_i))) <= Data_i;
--  			end if;
------ pragma translate_off
----			if not is_x(RdAddress_i) then
------ pragma translate_on
----	      Data_o <= clut(to_integer(unsigned(RdAddress_i)));
------ pragma translate_off
----      else
----        Data_o <= (others =>'-');
----			end if;
------ pragma translate_on
--  	  end if;
--		end if;
--	end process;
   
   process (clk_i)
   begin
      if clk_i'event and clk_i = '1' then
         if clk_en_i = '1' then
            if WE_i = '1' then
               clut(to_integer(unsigned(WrAddress_i))) <= Data_i;
            end if;
---- pragma translate_off
--          if not is_x(RdAddress_i) then
---- pragma translate_on
--             Data_o <= clut(to_integer(unsigned(RdAddress_i)));
---- pragma translate_off
--          else
--             Data_o <= (others =>'-');
--          end if;
---- pragma translate_on
         end if;
      end if;
   end process;
   
   process(clut,RdAddress1_i)
   begin
-- pragma translate_off
      if not is_x(RdAddress1_i) then
-- pragma translate_on
	      Data1_o <= clut(to_integer(unsigned(RdAddress1_i)));
-- pragma translate_off
      else
        Data1_o <= (others =>'-');
      end if;
-- pragma translate_on
  end process;
  
  process(clut,RdAddress2_i)
   begin
-- pragma translate_off
      if not is_x(RdAddress2_i) then
-- pragma translate_on
	      Data2_s <= clut(to_integer(unsigned(RdAddress2_i)));
-- pragma translate_off
      else
        Data2_s <= (others =>'-');
      end if;
-- pragma translate_on
  end process;
  
   --process (clk_i)
   --begin
   --   if clk_i'event and clk_i = '1' then
         Data2_o <= Data2_s;
   --   end if;
   --end process;
end rtl;
