--------------------------------------------------------------------------------
-- Project     : Single Chip NDR Computer
-- Module      : GDP 936X Display processor - Color Lookup Table
-- File        : GDP_clut.vhd
-- Description :
--------------------------------------------------------------------------------
-- Author       : Andreas Voggeneder
-- Organisation : FH-Hagenberg
-- Department   : Hardware/Software Systems Engineering
-- Language     : VHDL'87
--------------------------------------------------------------------------------
-- Copyright (c) 2007 by Andreas Voggeneder
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.DffGlobal.all;
use work.gdp_global.all;

entity gdp_clut_256 is
  port (
      reset_n_i    : in  std_ulogic;
      clk_i        : in  std_ulogic; 
      clk_en_i     : in  std_ulogic;
      WrAddress_i  : in  std_ulogic_vector(7 downto 0); 
      Data_i       : in  std_ulogic_vector(8 downto 0); 
      WE_i         : in  std_ulogic; 
      RdAddress_i  : in  std_ulogic_vector(7 downto 0); 
      Data_o       : out std_ulogic_vector(8 downto 0));
end gdp_clut_256;

architecture rtl of gdp_clut_256 is
  type CLUT_ARRAY_t is array(0 to 255) of std_ulogic_vector(8 downto 0);
  function reset_f return CLUT_ARRAY_t is
  begin
    -- 256 color ANSI palette rg. https://www.hackitu.de/termcolor256/
    -- Only colors 0 - 15 are different, and there are only 6 grey colors available
    return ("000000000",
            "111111111",
            "111111000",
            "000111000",
            "111000000",
            "000000111",
            "111000111",
            "000111111",
            "001001001",
            "100100100",
            "011011000",
            "000011000",
            "011000000",
            "000000011",
            "011000011",
            "000011011",
            "000000000",
            "000000001",
            "000000010",
            "000000011",
            "000000100",
            "000000101",
            "000001000",
            "000001001",
            "000001010",
            "000001011",
            "000001100",
            "000001101",
            "000010000",
            "000010001",
            "000010010",
            "000010011",
            "000010100",
            "000010101",
            "000011000",
            "000011001",
            "000011010",
            "000011011",
            "000011100",
            "000011101",
            "000100000",
            "000100001",
            "000100010",
            "000100011",
            "000100100",
            "000100101",
            "000101000",
            "000101001",
            "000101010",
            "000101011",
            "000101100",
            "000101101",
            "001000000",
            "001000001",
            "001000010",
            "001000011",
            "001000100",
            "001000101",
            "001001000",
            "001001001",
            "001001010",
            "001001011",
            "001001100",
            "001001101",
            "001010000",
            "001010001",
            "001010010",
            "001010011",
            "001010100",
            "001010101",
            "001011000",
            "001011001",
            "001011010",
            "001011011",
            "001011100",
            "001011101",
            "001100000",
            "001100001",
            "001100010",
            "001100011",
            "001100100",
            "001100101",
            "001101000",
            "001101001",
            "001101010",
            "001101011",
            "001101100",
            "001101101",
            "010000000",
            "010000001",
            "010000010",
            "010000011",
            "010000100",
            "010000101",
            "010001000",
            "010001001",
            "010001010",
            "010001011",
            "010001100",
            "010001101",
            "010010000",
            "010010001",
            "010010010",
            "010010011",
            "010010100",
            "010010101",
            "010011000",
            "010011001",
            "010011010",
            "010011011",
            "010011100",
            "010011101",
            "010100000",
            "010100001",
            "010100010",
            "010100011",
            "010100100",
            "010100101",
            "010101000",
            "010101001",
            "010101010",
            "010101011",
            "010101100",
            "010101101",
            "011000000",
            "011000001",
            "011000010",
            "011000011",
            "011000100",
            "011000101",
            "011001000",
            "011001001",
            "011001010",
            "011001011",
            "011001100",
            "011001101",
            "011010000",
            "011010001",
            "011010010",
            "011010011",
            "011010100",
            "011010101",
            "011011000",
            "011011001",
            "011011010",
            "011011011",
            "011011100",
            "011011101",
            "011100000",
            "011100001",
            "011100010",
            "011100011",
            "011100100",
            "011100101",
            "011101000",
            "011101001",
            "011101010",
            "011101011",
            "011101100",
            "011101101",
            "100000000",
            "100000001",
            "100000010",
            "100000011",
            "100000100",
            "100000101",
            "100001000",
            "100001001",
            "100001010",
            "100001011",
            "100001100",
            "100001101",
            "100010000",
            "100010001",
            "100010010",
            "100010011",
            "100010100",
            "100010101",
            "100011000",
            "100011001",
            "100011010",
            "100011011",
            "100011100",
            "100011101",
            "100100000",
            "100100001",
            "100100010",
            "100100011",
            "100100100",
            "100100101",
            "100101000",
            "100101001",
            "100101010",
            "100101011",
            "100101100",
            "100101101",
            "101000000",
            "101000001",
            "101000010",
            "101000011",
            "101000100",
            "101000101",
            "101001000",
            "101001001",
            "101001010",
            "101001011",
            "101001100",
            "101001101",
            "101010000",
            "101010001",
            "101010010",
            "101010011",
            "101010100",
            "101010101",
            "101011000",
            "101011001",
            "101011010",
            "101011011",
            "101011100",
            "101011101",
            "101100000",
            "101100001",
            "101100010",
            "101100011",
            "101100100",
            "101100101",
            "101101000",
            "101101001",
            "101101010",
            "101101011",
            "101101100",
            "101101101",
            "001001001",
            "001001001",
            "001001001",
            "001001001",
            "010010010",
            "010010010",
            "010010010",
            "010010010",
            "011011011",
            "011011011",
            "011011011",
            "011011011",
            "100100100",
            "100100100",
            "100100100",
            "100100100",
            "101101101",
            "101101101",
            "101101101",
            "101101101",
            "110110110",
            "110110110",
            "110110110",
            "110110110");
  end;
  signal clut : CLUT_ARRAY_t:= reset_f;

begin
--  process (reset_n_i,clk_i)
--	begin
--  	if reset_n_i = ResetActive_c then
--      clut <= reset_f;
--		elsif clk_i'event and clk_i = '1' then
--		  if clk_en_i = '1' then
--  			if WE_i = '1' then
--  				clut(to_integer(unsigned(WrAddress_i))) <= Data_i;
--  			end if;
------ pragma translate_off
----			if not is_x(RdAddress_i) then
------ pragma translate_on
----	      Data_o <= clut(to_integer(unsigned(RdAddress_i)));
------ pragma translate_off
----      else
----        Data_o <= (others =>'-');
----			end if;
------ pragma translate_on
--  	  end if;
--		end if;
--	end process;
   
   process (clk_i)
   begin
      if clk_i'event and clk_i = '1' then
         if clk_en_i = '1' then
            if WE_i = '1' then
               clut(to_integer(unsigned(WrAddress_i))) <= Data_i;
            end if;
---- pragma translate_off
--          if not is_x(RdAddress_i) then
---- pragma translate_on
--             Data_o <= clut(to_integer(unsigned(RdAddress_i)));
---- pragma translate_off
--          else
--             Data_o <= (others =>'-');
--          end if;
---- pragma translate_on
         end if;
      end if;
   end process;
   
   process(clut,RdAddress_i)
   begin
-- pragma translate_off
      if not is_x(RdAddress_i) then
-- pragma translate_on
	      Data_o <= clut(to_integer(unsigned(RdAddress_i)));
-- pragma translate_off
      else
        Data_o <= (others =>'-');
      end if;
-- pragma translate_on
  end process;
end rtl;
