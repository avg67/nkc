--
--Written by GowinSynthesis
--Tool Version "V1.9.10 (64-bit)"
--Wed Sep  4 18:15:42 2024

--Source file index table:
--file0 "\C:/working/_Tang_nano/gdp_fpga/VHDL/GDP936X/vhdl/rtl/FPGA/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\C:/working/_Tang_nano/gdp_fpga/VHDL/GDP936X/vhdl/rtl/FPGA/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
kJswNv5CyMI/ljX2grQDmLuJr7uKlop/E8q6ctap9pesVpBwy0jS1v/78wWusjV7gWqg7UMQZt9y
Zv+YUWB7Otn/iVrTEcXVS/Bvpps2hksuwMth2tfXoUB31IIY3ppCf81X4yVlUf79aJmOObVX8gHf
EegG450qoj3X9GgKN3sgnB5HKlY2Ey2FXhqRwXJk06hMnmD7gejY0Fg8Dd6h4GlKYxw+AkTH8A8E
hjngJJwk84crFuj0w3k2sMwZOwluqVM40n/xDBc4wSTsHR31Gte7Calg6H7Stj0O5pigFIV9WDV5
7OXHqTI0YTcMAamN/ShLDI6LKXp6yVollmnXcg==

`protect encoding=(enctype="base64", line_length=76, bytes=11648)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
rDOM6Qe+WHfCnM4lxqW1rlHMLvDkkDyK0bFW89bWy7D0LfRF9PDzvYN3FlYX8hk9+pTaxsLRaEyo
3Fxy95WYAV6qnDAwkMcvHtF3CDhfTqUsLVvZ/Le/k82/YwdmURA0YomoHzKW6S9jGJHYwUDyMk9d
tl0fKCd10BFyKMKdjj0qGWaLKpGLGi80zPAbDjz9D0ie0QhUPTTV9k3xhsEtvhMCtAVQJYChBucJ
ok8jc8iMk2zdrJHDWRRy4dABrKAIdUNhoGvzDNZx2elcxPTFaNm+1qNwLlqAIhNXlSPZj9blNawO
oYGwFc3KgVrnAofJTbZZOBhYKx56+JgU6+dXdaY/xqyPQgmxHfAiEI4hV0xYvudmYj2x8vucsBgd
5ePGQIkerzt5j59zfvHvPirWEtbtvpzbGq6cjIjjloYri+R3fxsp5em9VrB1almgn8eryP0ILn3W
nXZdUheXxmDEVGEAbN0IG+pFhFTtreirz7ZIYhW+IF9VzT+QPVsBVjg0Ow4ZwNHwdE1clqVC7Bmz
STfMa882+wCh2etP+tTwb+1YXYRAyShdXAhz0W1YX/orkroz8YRq2iLomD88nFVUXQf1ZEHQ/Hg4
eW+RPmHlT4S4pncrjBPxSa1BizMBBxTxeE65rRUlO7C8hluQAl9AxI9ulBMD5LD5wdHwtjC4kOkW
WjTgJgfq3v+L/IkoLG22fqh7UJHzBpTAH971uLmrTEaoQyJkP0SRR8lfPWJErheXu9yuZa9K02pu
UYjs3eZen5PgFV9asx8CPTK7AQj5T6eQQsNtboJcuhOX12lBLRCilXiUnD94OYtRKhbLrSddScan
UzF4Zp9q4M219LgKXnWPtdScmyp+RZq+dSak9ecoMKhVJ1teMSDT2dStBLAceTptBiUu3mPPWKdD
/UxbjSPFGnRI4FsY+N+9KVew7kBAANpprozFnEWfuketgtXLSbaghJx7zHe2bm6/V2YN5rZYo94h
wQEsUvK+GGMPvo+GHTNPWWhtpzAhhXAhdpQIJflG+47x/UkuShVLfE50bsZhEdAJQg2S1uEUvBOf
NVMOkKBWSVY9+RUkNy0iPjNpmCrh7CtJKDX35rMHp1cu3O67LJI9vDQsMZ0TkJlb211fRHj9p5HX
EgE32J4lZ/9miUg48l2S57JfmzeHUlxSaNo4bMkFPX86UOijrnQfTMfgAn8l6XFy8PSiHF98qk5e
dihpVQQPwdWyEAQGLIUqU2oVjs9fxcsr85Udhg1Exgl57EEbft73v1Lbu7fUI+LDpmWWzO5NOGjx
q9zRwsAXnFwku0cUYtWBAUdFvdDhE1/08rF3oCPxsyJ0Fe+JKv1KoGNdWmYoqFskOh0lazgVG/wn
All0ojYGEb69opC5JPj6EsmFkMD0ZYaGic/eVFHetxtkDDNyWV9DVvZIPzd4K3PZeV6F4UBcNbfl
yjgz4Wz6Oh2NIJ8uYjqsyeMNhmLjj1igfiktzw73eOdpmEaypK6EVnv0RQchyoVliKpp2pBGd9Wc
OqE48dNvDtpGUKFT0NTtoxDTXZL/GbaqoxK2vT9IxqoODPy7uFmpIT2u5mBtVfrSk4ZTlDykiQF+
ABcvOIhWQ9y1p5mp2+MO7IKwCRi+0PbfKsHHyrI6/iC6nT98UqpZcYyu1pDFbeNgRHT/ipIt5zXp
uFGUb9Tcq6FmTGXcLpGSBFAvwKnwMoqmwWgWO4ZD/fxgum26+JY2qC4l7dN84Eck6lFnGhquGsn7
vhRheViwJG+5FDT+gKsBdUTmoigyIwUq6CUPvpJCEgPcK0EJXplzFrWIct8eNplPby3i0bY6wqxO
5vR15fUK0f/McTOU/ERlTaYs8HI3N1lV/GW/4L5Qot3LheOCHGd0hEg/PHAiirzLDtu5X0oosFsj
REn83nUU3YgaXtrM3yE4ThTpR0FUJx8CMvHu36tr6tSoAyZOPy9dO9cmTi9yCVVduYl3GpzbrK1c
IoAPB+P4/afyqAdLSs0GEGtxidDrLx8Pd7kqvitIFasw8CRmbQsLnhldZrfScuxv+ihkFvd/i4sR
p4up8Nkc4Z24SN7tE3T9kByBtDxVpbw9OynIKcjRKa2gVx4OfFoguNtFZivleFDNRd3zn+1L198d
rTStXODERgT48UmnQmXn0yRhrbJz21ebl8AnEPUOBd8mGDb0BqHJ4Uz8UHJMbhyt1lc8g8O3QK0b
ziBiDFp1uSpA+DG9+3bb+NHL3AXSHQTFgfoPRBtC+Gosx61EUQDalFdoXNadgGHMeKWQl5vqALrI
gdnsemTfihfq/8PpBdDeI5CD2JHJ5f2quRaRXO11skFOjASORSK09Qyk4UDi2oLIXXIjm5OH/WfJ
iK4tiGOty5ewXwFEHLpPo/yWuWWNC2mXYTTkYqbz/GHr8L/MyEy4TlAOh4PwX6rkYU82j230Sw9+
D4q2X6sKoXf6uYU2J4C63QrdEs7TULCtr3JvXl/mev/3tSX2f4NwLshckhc6QJWSrWXsm9u3mEle
stWD2mFQBFO8omERbOFTYImWsndkXjHpHyQjHC1cMxubSxofuiYFF0/wyH6VUUhHC2sKiHMCr1xY
aDgf+0aYjI3CqUws3d7Gr40eAIwuKeHD3LIxTxKlx44yDKj4GV7AV0DFHOBQqlOxFXez695p7w/J
zAuZTEuboDHqW0mhfB3D4OcfuJBGEKlFFUxb+DD85ZjvaiDsTFrwnc4gtdJkMqL94PjeweBp/4h5
GHF4tSpukexx49wFHCU/jIS+3tbR9Fg/NE2mXvmP1DEydjZMJV70uyNs9yLfM6jUUvpG0hmBSDWP
wwbuW9ZZguf/N3HSfvHm9PlfFIx/u0BCBzX9xkH0QGbR2e1M4qUTvVLYivwX7mUfZHyMBNOUlJRm
SKIPlHsNE7QmFhFQTWV4bKaUWZUsm0r1eHUY2D+USFOaMAvqoCHQ68gXqMywAqiZi0hAEaIr8Myc
ajFAx8M/XMcIogq78p3Gw67c94c2hg0vUHpO27EvI3kcGOzbSX1A5xUAVpsQHWc66baN7W9ASi4B
9yW4oH4vDlSBhdq1u5HllCFmhFv5Zj1xipL/2xbmp7BzBeYmKDCDEHMYFr24Z2eZuJdMlu7vv24D
5XZhZGPvxujkWyeVUyugNyGV9R0okbNYbkdHW+jfRheBK7Wn+Jsc5NTF2jAAs8yWK0zZjswwxW8C
pB01NIOVRjGIUtpq5XvdN2EhWIkJ30ZS/YBN1IcEdlU6iFXAfZzhTcmwjjkt9xB5arZn5QZVD79G
Y78lEq8Sc0Zi/zrBWuz/kB/LFbJccGa0lolQmSsW5pltAro8iCD82Pvqz+Wcmo2F34/YAp3iKFjW
VksWvMHkcKAA228cTWaae56woJs4L9pHIkNi+8KgqlJmp10cJsnRsL4Fsp9y0quM5qz8ek1/CWnH
fbq0lIP6inLCvGJM9z4O8bG2thWxpTBBG3Oau5dDJUv+jUx23XEqZBi+q1KmX7oR+maN7vHZPoPu
mqi49fGJCFQ2bkULM2kolJsRbPxK02W+b0I/0YUPGorE6v2ubbAtaNE7VCS/RxraHy4VqICHR9bT
8kixTyg8w7v2nY9s802huCc3wsBo38GvJcKN9u1yGyCkKWbuzzMWKvp+HBolSOAWBzrvfnWM0tF/
2H1vALZaQUjWw5FHzM/0lLF3+pV2WcMDOa77d9esQncDEXAwXSqKBoYiv6hLiUKxwF/n7wkuGkba
EGV4GeJVHa1tLuIPeeT+iZ/aZ5bDUp+0vfy1L4tBip4haS9OzPn3TwEGAEwcPocWXkSiRDGaV8AO
bhwkt04iniG4OCUBoulslpChCL1/pWeycm9++lLF/JjqnzyGrtqgQ2HgWwEOZGAlal0f98l7m3vg
i6XqD3bbFTGUZZodQqSGNaqib9C6XZrW5NO4XcTHakmSbwU60As+9091dNo82dugNZJu0N2sth+a
Lz0TgcEiwla6PTqeVmxVn8OP6fAdClECskyFBuQCxu5sxHpVw0Wh7/MKwUpqq3Hs7Cv1TnR/eHGW
Bq42b/Aa8wH0aTDj6vBARmf0nb/0a5kdG1gQB1EB+l2ViyPckzlWLiDLTxUDxyEFfK1xXIgJ5wm1
SPqT757TQa2qdMmzYJpULljTBKwADYOBA38BEQP2EWY5iDuMw1EgctOvk5V9bYpehlubCMxHfsL+
+KvbqsZcrzCCakstp4zbZEDyP2XO6+Rw3ZEBaYoKZOgR2D6wMv91qkiAqGxHUtdWgS66Kf24xWXQ
CO8g2yhJa9Zhtc1umKth73WiDWHzqwFUrXzptkuvVTEh1yD2Rx4nEe2IM0q2KHq7fwCotDYKa1g4
bqXiJFZcDdiASEOOo/fRTViwAgrc0tjP9YDAf6NMqHiPAZss2R4hlsx37ep0kSzkpcyJnlwdybHl
bzN56VR2VIL7yqlrWlPISqpI6lPFIA9rabwlb64teZZ/AjgVVn0TD9bnamHXxK/MSetQdwa8DG6x
7Nq30aLhZOgK+yUUxYA/GV9uApF77UKWlJZJVMSIMMyDOgbuEK+YzKSptJ4GWPoSUhO65q1UxCS6
lV4JFJivOcbAy/mCoZnCxmLBYL+/f+73aWjZogj6I6+rtQnDVufBlQvsSXguz1I/dW6RdTl9fpwa
AifKowt95gUeGsR0x5fIzWYJOzbiRdvg4J4SxF6gFT5hi5QOHCRDLidRYlG3ME7oKD5iI9T1pygk
t2uiluIPVq4Rgv43N0emMXoqI+16csBGhAbF274leywip30j8qI9ItMZVp7kT1b9BPvSyA1LqU4Y
O7OlisF/wJj2V3bRvhTxV2bQsMrTy+fdOfCRRQ7Rty0Fct7p/XR1gCfYYP3RPA7fLp9cSxg/7GJ0
3DYkxJeRJAJEyrxVkwj0BZ7TngBVzID5TUUeR5Mmnbk9McW13y6Wp4ZTysvQI1iFVK9QKIjcdk9y
pt0noOsyM1XIoxEDePcPx7SmHQh0HbtHPV8rh820+MrdEBvH4vc6WB+7mzudbBzrPxbPAv50NMGe
YcA3lk8+oJVokpwYQfD7OAWhpGkLh8b++IwxQNq+WXXfmIxIlmC+OhyCp/WXYjsZGNJjtciDOKbz
ApOlqr6aojplLaGu2nPC0LAUflTW7QH7LKZ+VhYlr2I/XmjNRYdh1A9eXqt2uqW6eYvDutzfaCdC
zmy46MpbW/BcBjCqYuBvZb9WgH9DCMvRf5fazT7L0NqYwklwHP6Hz6aCzQXqq0TYiHDHrRwiwWLY
D//FW3Gl5QPxwTVd7E7SVyegSYjNlNHBVGfJJFEsjDg0ClkAbBszoYr54VYfHPAkIVjAag+PBW05
0awxRHsF4yMXEo4wd04lwLLebQiSTocOA7AXj0Mc3kWeX3QxNJh9/SGqeuve6yeyWCCrt+uvs3BO
QL3hRtg3SLUNNTbD9bCo7mMDqEqFtoyrP0NYLizecQ+ZUQ5OOV/TuJ2l4IaL5zZHO8QlZqUFmzdq
Hm3zplErkctPGSPrtOMsUNsNPyJoeGcZZ/HMB2jmETaT49iwKibTAKrjAtI4YHgvvnDCxjkx0uT9
Jv/2s7xwNu+amjYLoLA3mE9tE5OCwRe7SZMT4iYgMqerT7780ls8KI56a0Ag3wY/yVRSm4WbzRFH
GO4ReN5V0U+zkYFN3LrQdeoEtfsfhtQmpuwDm7PfrE8iGR0NX4OdxuiVv0BlWkVpZRtY7cMXwZkl
EvpJ9jY4Ph8OdDOuzYuAMU4q5t3Xi8ij38FR4kIffwQdYjFrnxnxLzZlq5bN3CaQKl5u2G9OJbwv
R1w+CQZKIgDQPoFd9jnYYVEbh4GL7jAWldiMhi+S++Vun//T2f6g4mvrW1Vkbs+q2ShAdUd2hz5X
ir01zSYJD9f/LnqEhP1U3+qNF1FVtLSZAFfWApZmMyjZ9kWY0BfOLqo00GZCKV7qcX/AEeJrhMft
hJ305XRHHoXLddB6igdxvMWfQ9VYs70w9BwwapXTGe6FEPPL8TwQkTP2qZTLGE4Y+NKl8YUFVmqv
1t9AiOTT/CJQcDxSY7B629VaXq2+iEcC24ydm1+2pgw8sAZdebl6HWPCse4SX4sEovXSLTgj5K3K
uYa8V9IMwGtNunYLDEVZuVq0qYOuErMQvDgH8PmnTnMT7XXnf4uzRB7CiKDnhotoHKcBcCSn7Ymd
N3Wl/NRNz0KW3KBKEdqOcnozSL9K42Ia0TtqQMCdqf6HLz1PZmgpU2TqDgo6SWODkxtpgELLWjrj
ut8UdJYQO2V0sSdunMuZyf8nXCpnG4Utog0227l6NgVtA9aWDRwhzA8kxpuYzndkxHWV+9tMk9Ai
55Ciy2g/0NQFs+0LyoI87peFaXqdqbavYOiT8fgT3bi3uC2XDjjlIZ41OvCNk35AzMb9m5N6hWU+
RYPNcc6OarallmxusxkiyvUTjtbDQFk/4XktHzzib2qavYLwKsz479Brob/sWndG48S9TKWAJNVC
9J849ZyBxDOJ0FLZkiWBD2WkqfdDv9xwEY10ZI3xgOD1+MwQF6ttWOSH3xW8GtXJnGURFdKxOOt3
sYwzfo2mdn1FkWpc3ePu9ONy2CQgzdHbmm1rYvgV7awnVTX2XwtzPOcmCCKBT6fy7CfNKs4ntFRR
T9osEKVVzAODZG1RnXuqKCazyl7oKCq9J+bW6eqGxuTnyZZrK1xzhHRU5zeDrJGZHNNNQVRpe5Tn
hQTqHLULE5jBeg/D29mjMVB3oojxYIxtwR090kLJG2Cmt/Go/6KF4l/7NWu2AObvgJhEyk2H0n84
zebhXccELcVJCpqiFFy1JvC6/9Rs6wtqOnx0w4AgALk8E7FHa6yt6xH3jQ295cIoAbiuLHSuthsB
zlCg/+IQpMmUxqa1rdeT5uemx5MRtmEm+3U9hLILDDBBMAyPZQpvUN11crWHidsNdP8FOB8ZSUR8
83Xq/ud1pSS5dz1f+fhjbPVXPEwo2KESgU8egnqyIssb3otcDiCMZhb1h2/lRRKbvg+DnpYZJ3XP
qX+FjlvWhN2870LJTjyhvnjVJC2kDrQQh6I43CBoHB2Nve8WL+ITBKnHhL8VVjUHVr5G5+oI4/2x
J24xkqJICp0ljoWTStRcQe2uieYcu2tLetwBPo1gvbvGUnc+YJzVuVeuF+4lHbgUc6IyX58VNSVi
j/cCixpWE38DHkFhUoXQSfC5bmpQbpkTnY4DVJY7jbrDEZSuM6WpkYBdDjKuMAQ/Kx1JsseF5cW3
n6O/01g+RpJY2MX/POVe6Qeck1kohb29y7sKe0f5CVThwQH5JQW4vKMVjPkT9tMbpQ4Wn1yG3PK4
mVcPcrLdrO9VzBIVp6akXjDkDRPZVUW9AYZLtqAqDHUh2J4fFfW+vXNFcjhFb+8K/o5/XZdCmMwc
QIWctgkXp36SDGJa9R1R35ZPWQkSonzm/2xVmsU5HZW+ClyLrfKCIDFSBNkockSvs74656ckm9Dw
22rKDCKxuFRdmmcYNroqh8yEWvJ1clE07RoLZ11Y53Pi9FZGksadGQu7IM6xwsUDNeO6nXcJ2/K5
W01sbAx2mE1PEsIsHCZRvuPH8ur2sEQzAZt4rBCWk0HRvLzCJkSvYel0fMUEP7LQECUju3BxSk06
gBFqS3W+X3vffnW+6mgajo8HNkyWFCibnBQOb+EjHv0YPQ0aqSnXQSJ/8A5uRwDauoTtnQCo7NVD
EB3r743ueXamXuQiMpODkuCLJcqM+U4qohw+BW8U3bJHkA5HgtWRAXljCevOxSUFdZK2tj7jrcj+
UwntCuopxq36p9V4r8YhevWGsIESn0KKdJMV2P+8ioSRe0/uLmg6sF1xLFkSZMy88stT3vDSOxNi
yIVoPeeE1HGCyWCOAB3tM+5Kp4aB8TBaFQswOzfPJ1d3+9+OJvHgd/sT80SSP/BWJhKTBHoKweMh
+AlJKcFmQvg+/sRzk4IwSpq/CEfis49JvXECrEUCgWz2KkoF4RKmmtd2UA7arYQGxY9dtoM8SUvR
sI2C8Ao0P5Dq0ft/eJVc7eMy9KybL3g/BcFpjw1OZzd70chj0sVqQEIvDD7UeVXznPCkhCkdjMAJ
NWJTVAE3wlgapWxD01nnuT/VsCb2pCIIA/EKJ+VQtXgRmZrESn2IHlketzFFAStNqAlWSiSsRn0v
CyrL3saEu1sqQJxXYOSs0KJz2e0PS8ubMyG4n7+7gg7HMaPqyJWJ+ajrMuZi4STq+et3NA1NzxBe
RvaQu3mh0myBFIPNvgBVZVxxViKEFVOzVeYceXXW5rfxXrQoSiSWFTTV8EDLQYx8OZItCGkIFeTa
P3iodY2aw+DNdpxqW/PearFWFMfpBwlXXS+fnphKq0W8lxfjpJakhjTGM0Q+FjONK23KqU/O8Cus
n8DjuXqtEA1kKz8YSuuZPQUXNHI1qCaBhMsjGjHnqYG3255UAv1n2T455H18m2nxY6lNSvRtx8+P
VxRnX1f4NiFniTeAeBXZ7fpp3poSHjHViMMwDUYwMtSfQOvujOnpYwquTVvN6xykmE32xLNl/RlX
Itnb37QyT2jj7U+xiRfmyESgk+DNIslfiAbCrc/UxwiUEtf8N072VMEM1jcli+CLVPjCi+Lsw8bZ
bvVDcAvA6lkrEG0WPDC5OuicYkj0I5HWDTeK0RFQBfYj2NzE53E8fGLGYBaIju/ktaAVIS8WgpY4
NxLAzPfxVRxruVEpXJfq5V81QMDjD44r7defO5InQRQwlwDUXEkpZ8mY4unmDdcfr5ZM/63vYtcl
xxemCbYDJOlsE99EhiqrTlI0R5dfwxjL0DfdeAW6SP8hYoWR3CGSBAAlOEWmc6ERNS/fhmuUJUHk
FJgK9SQkHrDe3mXJt4sZwv6jBdC2JrfP8ucjiM98i3RWuPzeXUltfASlL01AkL16Ap6t9YMnDPLZ
EKfX1PmYhj7bbXG2GjShZ5KEg/x4je6ewNX+JArSzZi3SpbfnUm6EVIog24pe9fwZq1JHSr178t5
VeqMNtSOwv7v0VYjOP49tio2b+t3wqXGMmQBZBZHwAFRcyQeFRMrEqKwBPM6TzEmb6Jsz8shBRAM
IkeH8Qv8YS7nHF/R2CH4G0wY8inndZBO71WBI1ZEKlm3++w+buFOW/MIoHwVZvpIrjOPuQYSAm5o
SZf8mN2r18dGrixH/6lNaAe9Cav9W0Z13msIrwAaphffExeESd1QTOpbrmTYX1418c2JMRF2Npvj
1R/U9F7xfdekutNEgwhMJmZmEcesc7/sPZA0yFCPTNqBhRuwc0gJD5dgbqMClx7ET9vF0jeMfoXP
AODYIBiuFbfF3rjyz2TTKx7/QiqaH1SC5zg+9W5as14dDPkI4hk0bo0M1cXfNE3rjmo5kja1CMTP
lCoeR5RafwkUudD120n+A3JRL30hUnEu2KELo9K8LFgdzNOPBtQOKFJd7JIwCEYUQqkr5zA5g2Mu
9XYhbHLa7cq3kMzOX01vM5sZUjXVVJoV4bTSZ9XACbjTIuGc/3G/8jdCLJjUIaiFyWyz2h6CCWM5
b7EmoIRQpA28BNcCRRkYwXOmByDLvhUKZ80AgWUXm27XH6lBWsFjvgAiTKiPnGBK7NUis/f+Brb0
b/zWLVJMICGW40eY+4feHXFMWIVqApKR2A1+IuHmFSJoHoGXw6Y0pyjFA8uagM/+fodTLtHeq0Pm
SlzORsC1OoPBwCKZw85Xb/yeyiBNEZiLBNgr5TiqYjwhzhRMJox5kdjveO1W/DCNd+/SNYELZ9Dr
qz8EWGlUT4JJjxdNmo23UQlxHIF0o381IlOvA4NwTOkE2EFUIGUVFbAYn4G36x8ehcSb1yaOQPNK
hiQZM4kgQywuFfgU75DlQrbEJxoR+ShNS7bG1jowbGCC5iyxuNLc9++OcY68eJGNLxYC5LuDuTw8
PgBtHlnZkO6c1JkenXyTSX+hwtdtrjX4gsXvigsGfukoOvzymPNZqTdj9DXqxguCk+cEKbe63A4c
f59/b+c1r/oOXAU3bZkrEeNQktFLCgs/SD4ImXoxLILvMNgUdikaxUdQCssQ/duH9g6ubklPONvV
vLRcm6kNyuJqS7GQ13r6SSpmcsCdsWSNS+WVvm89PuaArnav5qrVteNRTpgP0ZXxLOK5Y3ySHjF2
FNJDbZubfWz+ZIxKvXR/6lirIiJg9bkF11fVOumSQg8CHlDZNBqO1liHY2K8S3KSFKFJ2IKmUUR+
rYQoLfgP3LlvQYea6iT3zFl7rrK/bMCBl3gIWfeQbo/3s3myLSOLUSW0jlUpQ8oaENw7MtrcxlFD
al7ucJBROggQ9hTF38uZB96fEMbqqRAxRMWYLuqPaeeNA8Y3MpUAQ48Ush87rNUnwWtO+MokPZqx
9q8qzTFBlMz/xazNhSTog1/jhnwHaLi9H9afbfvkQ+WLlRASmaTy83oxIA3O2fY4XvBfhefmHy5I
0WVcnWW6Y2hbv9L/oiW/TIHV2yxcgr7UMyn8gr76Rpjlnc6JqQCythiFsjidKPFwbWYAD9ChrirL
+jqwZDVqf7oIPNutWpUMRExSgoA5syciXiD7tiPC8T1BHgdOZ8Cu8J5CZR8rj0iZ4awyQDB3HYuy
gLK27siy3wk2j01KkimUzU/CG6y3r9//eg2rAskxkG9w/zIlUsF8O/YM/72YFmIjgwUIRIxkKY+5
i1ylVaIXi7pwMq5ZDh/Wp6rfY4XbFcy0D9kb+tGaKnjgxBu6PKwMGT8Uy95Yj95JH1HFfCHulObN
Uy1rCZQPPRJcNXMRNaPA7EO0lghXHGv0Yq5iF78GiCidwoFT7Dcid82S7Xe4WLHpb/p7XuXABVks
ZZNNK/nrq/XqnBJkqMdSFvkqVK1yppyg6pEMJvjLFI3XhIY3mpPpoVzSmAsZ77nlreQ4WBt720q9
/kRsQuKj4/AlTr0rz9BulrZiPB+dwPUupTgzm2IKSvtAWiN0/E5c39RplTg7lCx/nu1tXEfLCRmH
DCdLus6hFBHrMzKV8Whl4qV7dlu9nixghE8qbtliWYfz9APuMKnkjx2mVRL/1lE0JcjjaQ17A3wL
jt9zx4liEDhiB0EUUsxTox5y0ONKdzNfoCIBqzsufG0rfZET3aFKmA9qW7g59YzKbTt2xcqHm/FL
BzDjl/RpxIJ7WH7KGNVsTcn/5DLXccIILovQUrShnhHszuDvIOYEIBYoHmafroF/9Rp1qzPQBWGD
xOYXwm9dcDRviwB3i82fqRDrB/baCT9XoOpu4GaaCU3kFeYUeCurrIMNiljxqZetk21N+XJQ/5yR
EGQ2zMUydv3H9Gl/zXlQ5B+vKHDFxGVja8narizGbboHqyUGtdFHJoY+dN1gFXLAqeXfqtvrsLGD
jS/d/blyupOpp8mBKFBab7yyla0Inun+3KhTESwpQ6FfE394lZjj/vSA8D0xFB7bcevbwN/OMRzh
FXISEj0Bef5rytJPAPQ64IdfhSHBgCz0f4Pp2j84Js7uU2ZFMdXE6RgU/5tLSnB3TVUoamqOCIJe
wJntkdJTDMjAAjCM8Sd6YTj6Cmhcts40VbI+jt6NCQNS0lLqNwmIoQVP4k9Crrr7kF54m2VLB1jS
D/zudn7n5UU5JRwWD4fuLxclvcH7YTivyjhS6tZ61oXmC3yx9lJOyxjTYt8cdF6TZK4+qpcFH8jN
mYtfaQwdwW07ilQdhhkc9h3J7S2Y7vEqCTqTaHntJvRcmi/7NhA/vRi9/wQDWNLtg6wIzjD/J+l7
+2MrBVpCFqWLpeqA11xS/b/CY8ZodH47ps86BUPnQMeF7uMZIq1uTrTpe88GnZ09LX8Z+7t4UJbK
9B7xE4OAUBHpvch7PZntPmPsz7BqOI48BRKlWIcB+Z4m5/RZ8JHR6shbdR/TAqxn+1HATNPMXY/6
6+ur1jbKyzXVAf9xFYJsWgplj5sE14sgGtLet7kFlAreGyvjf0QE5T03FjYzy2yNIJRsviFVfrfV
+yTeBcdBcbufxUr8j8UNdZ9HRGc5eBip1Tr3/Kv7FlkuwG1W+fGg66djApdYrgy8ZFO+T6Ev6PRL
NwDCGnU80fz07ov2uIMeuYPAsdjoe52FHPxlift2q8k748o2hjItrBAiaaE3FtC2W8Nfsr9/WEW3
baMFOmOJ4NGun23oBky5qzjNtugycGkpnGo1pXPBDCzZZ1jsq0DF3HfQRfpgbN1shd2r4kurSRhr
Jto//WHtpJJDZHREtiRIjqNoPAWb/Xgty++tZNzukA8YVUznNbYayjmzaZF94AYxUvCDNHtK5mEt
UBuPhMDHKc4WZccJf5IhjiIr7fzFQ7X+tpkTOS83Gvet4j93lCYl6rmxMWSPxGdjh7ADjIeX/2c0
Pk3zXOjmBPy2bgnfGrTchu98CLXPhQGWu2qAk3GwSDpQ7PeecIlHQ6JL2Pw2nt/8TFl+Qw/ytTcR
GE8T6mfL5Vv+2xpp3sr4t99uiZhz+wJpwstFkkjxYJEpuFuq3UWPrUtIEd+3qCo1qpKExgDG3a11
919jLvkPVRMV8R4+rJ6DpCIzoAJLTSwmgln13FksPxMqwtppOOiF0dvMiq8MfAL5ICoKEaQ3rh7k
n4ZISXFAIXrArwanWctbpg23DkNb7brFsLi5SONVD4smJEvifZ0QvZNzfKS3YYGAmErNZjAYDgxB
dTyjVmqp0SUFHD1hsLNzlAi/Pg2a84db6AQuP5K6ops1bC1NJE+CHqAShD4txn7zU9DnMA2myStY
J3z6OaAcMoMl/o+HEFyj8h7OYu8x7o1FqHGYlpCBtZrcAyljXKJfJ+QsXAOjvhbm3/ZmDoY5e6vI
0HemOJremObhd/w9gfK2QZ2iNt+fhcrY2b3ajyPQcU4oa5C1HGuk+ZQGZtsNa21w8aDtSEbCSGek
8o/xEuiJl7aXgVN63INQbXYmJE/K0rcX//g2T/QW4awy3z/VZjGJN7a6Ue7/QJryV6vDLrFbRcIr
gRs/kGMTAPDmgwMuAVAPCKHNktPizvIH8pUPd2aKoEOFTWFzyNtGy/kR3HdaxDnlaISVWbSdUKYT
ZJVXX+LFYpbU9w69Al00sYdWX2P8SKRlpfSjxMbpXTXhUVY8svz6ao+BkIfG7874372f2N9z8esK
5Sx54S1HivhxahxloAI458sL0im9Ssq5IFPFG0C6Rm4eB1V0ztkGrEIFng/ysij37AK6hFfr+7Ag
yP5K5JBOA+UqBCIUNZIgEc5OXwqrbYj3yWqOs2SSGP0El0bkaMoZxMxcr4Mqt9+o4SrxGQRuW5UP
7q8gbUbpTjkzsCNPOBXm2A8hDQgANZAb3y3uIMbcK49QQ4dNu0OTaWHr0pTreOI7R4GWFBWnP+MH
JXJFhgSCqqu+w9dw4MKqRHwm0sorwGZ1NwG2ZubOSUfCbhj42JYDdSvbGw7Y0yCC1xht+4lJLvFT
Pz1+kfAVucJOF63jGDpl6/dGcsEErNhBfJK9Y4hgxopsQUuQkWfJh0UmvuYKz0X8BVg/rjLeO/ns
yE10prsi5CzMcJG+m+WLMbUZa4Q/nP0aiujNX7Qzrlk2PWZt/BMdeaDuEBYaD2wemSv23q0tO7gl
Mv6kAVesXDTxrGMlbXB9cwrpjMw7J0AOmnsev2+y6GWsIT7SEKRFr4hXnnIPSSim1esTg1AVODUv
2ppaWNOGLLW43WBiWieuxXyCICYu/xP1NObd8+ZDdmGJGvh5/XiyWYraZsszj4dbK+HyTalq6VLE
JKt4LgQ9cluOp/ZyuE4LLCnAgpZsMhQTNEtxQ++ZLt+EjYMVvVrSyX7OMhPPAQIsyEw+Kqoy3WMO
uOlsLTD+Gafll2sPnTbloCxALJJh5FZUsLwL2eGE6IBAeXgwAZ2MPbieICvukASdKhjvirDLCuAf
obHeZ8T4qokziq2mKc5B6DLnVwvObbDIXjzRUGUsRGThsyn+PV0I8dz1oH1OFaxHLeb0zmspA38G
/ifzP2K+1FMVG11B9qBsesy6zsdJpbat+konZhKuOLBcKDLW0k6y6cjZqNdinVKPK3u8bSlg4tsP
PPNQBgYuYXQsqoR2tk3LWK7nN3r+rkTainWDeJdUxLn5wI0UlnQcy+SIA+Z1JUOeEBhWvoMTD6nT
OqbeDnLeWdr12xMQ8gqj5STGnnQe7xLd8eaJ35TEwXw2EHeF30iZCKQAjcmn5GUgWUqZitx2jtFN
pJ5f8zswAAnqiIWfvrEACKzgpk7Qh7o07yy2RtNUVaJME7zilKUlCfZ1jT9kfShdMg0ykdEuXbS7
6vHyY+nTOfLGhdUwxPGb/y10rKX7y2DgQ1wxuvxrAzlEKrOfLAj0D4KGIL7ydBJ9PclzMD2lyUVF
wDO9x71p1awfqLxoL/NWSxSfT7/VIons2vi9uNTVSHTnsGiMQ+V11S2OR+8d62egzcWgOF3exunp
nvIOaWTZFUdEXGI7Ar2fvZGAz4wXhFbeEAPp3k9940qrZtpIk2XpkFXS6ScpsiMVB5iYxyoEap7/
DdDyYjoGDjUkwt/AeL7NxKD5AnC4iEQjtaGsQ+u94Ae5aHDWT3mxvNXj2a/zN3tU21AMGGZRMyvy
ev4h/rgo9y3OD9LRVz1guscG2hDkyoXCbW1x77RTngzuZav8nD3eaOLJwWsUxy55F6MvQWZaz2T9
5SFYGjg2gr5MQcXgTYFDswWTUePb2BOW/xrRp/xVP4sm2CpKyzLAVyhNcue4l7WvHp6b6LWD7mC9
bfrjCrhuda2cpKe2gthgUP0LH059vggtAcV8YT1qHGT8kI9CJUxVQRJXF4TgeAh6azOE0qXBoGSK
/vgFB3LYOF97zHQP2UKYtkng46PXFAt7okB4zpVLdPRcMtur12WnGLPG5VabUn+4bYvOxDY7wK4H
0HKq0KY6ohdw+JwAOB4Xb07/ubFv4ux3Kr6CXFciogR7OHvvTS/eWH9p2ligRtWmJ9s4rZXum5zz
NamMo7kt6+Q7BQmS1MvEwaMWLKAouLpoFI+UQcKNRaTV8YS7AhGQ3vH48kSnWMXIP3o6TR0gTdc4
ikPaNTsg9MUieSbGDToRsum+Cz0GHBZPaI0VoRQ7mW5RYzUl0ZI753atQj58E86NCf0YVWUfiTvS
QEw9Cp5Ay0psvi6B92tFgCILT8iIShvAcaDdDD0Mhh7wujOpk5WUH2wlI0qJRcc6zBm2JM02aAYb
afj1o0WbIId17PCLB/17TIHdgj8kfeuktvUQAvNMx2rzEcT8Evjk5X4kwpgsBwO5dD/DvSikDxb7
qrh3BOFoaHFfm/cRS8EYUauQkoNw1VEmOAmYBGARzthleZU5gKjXWMlyylIleq81AxZqtFwIz4+1
U6vLF6f72hPJZjjrV7XeLwSAXqAUglIrnHkvoU892OMTABc/aDDqsHhFrHfCZeFYOMTiXeVSEoK5
Wqfcy56F35f0e6QN6xnLHOscSW5tIwsXa99YmgnbgL3RMWZ8KN1pIC6kUlaLmSTpdHKW8dhLU/a/
uQekwalZ3rh6wiIQBpxMa1S1fnO5ZXymRf954YZffEwu3CV2p2B6mHUSl82RVn9mzMeQIIqhpzbW
RfiOssEFXNAwsDiAYU2iczjUddc=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity video_fifo is
port(
  Data :  in std_logic_vector(31 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  AlmostEmptyTh :  in std_logic_vector(4 downto 0);
  Almost_Empty :  out std_logic;
  Q :  out std_logic_vector(31 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end video_fifo;
architecture beh of video_fifo is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
component \~fifo_sc_hs.video_fifo\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  RdEn: in std_logic;
  WrEn: in std_logic;
  AlmostEmptyTh : in std_logic_vector(4 downto 0);
  Data : in std_logic_vector(31 downto 0);
  Empty: out std_logic;
  Full: out std_logic;
  Almost_Empty: out std_logic;
  Q : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.video_fifo\
port map(
  Clk => Clk,
  Reset => Reset,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  RdEn => RdEn,
  WrEn => WrEn,
  AlmostEmptyTh(4 downto 0) => AlmostEmptyTh(4 downto 0),
  Data(31 downto 0) => Data(31 downto 0),
  Empty => NN,
  Full => Full,
  Almost_Empty => Almost_Empty,
  Q(31 downto 0) => Q(31 downto 0));
  Empty <= NN;
end beh;
